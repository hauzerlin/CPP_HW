module c4250 (N1,N2,N3,N6,N7,N17,N34,N51,N102,N119,N18,N36,N54,N108,N126,N19,N38,N57,N114,N133,N20,N40,N60,N120,N140,N21,N42,N63,N126,N147,N22,N44,N66,N132,N154,N23,N46,N69,N138,N161,N24,N48,N72,N144,N168,N25,N50,N75,N150,N175,N26,N52,N78,N156,N182,N27,N54,N81,N162,N189,N28,N56,N84,N168,N196,N29,N58,N87,N174,N203,N30,N60,N90,N180,N210,N31,N62,N93,N186,N217,N32,N64,N96,N192,N224,N33,N66,N99,N198,N231,N34,N68,N102,N204,N238,N35,N70,N105,N210,N245,N36,N72,N108,N216,N252,N37,N74,N111,N222,N259,N38,N76,N114,N228,N266,N39,N78,N117,N234,N273,N40,N80,N120,N240,N280,N41,N82,N123,N246,N287,N42,N84,N126,N252,N294,N43,N86,N129,N258,N301,N44,N88,N132,N264,N308,N45,N90,N135,N270,N315,N46,N92,N138,N276,N322,N47,N94,N141,N282,N329,N48,N96,N144,N288,N336,N49,N98,N147,N294,N343,N50,N100,N150,N300,N350,N51,N102,N153,N306,N357,N52,N104,N156,N312,N364,N53,N106,N159,N318,N371,N54,N108,N162,N324,N378,N55,N110,N165,N330,N385,N56,N112,N168,N336,N392,N57,N114,N171,N342,N399,N58,N116,N174,N348,N406,N59,N118,N177,N354,N413,N60,N120,N180,N360,N420,N61,N122,N183,N366,N427,N62,N124,N186,N372,N434,N63,N126,N189,N378,N441,N64,N128,N192,N384,N448,N65,N130,N195,N390,N455,N66,N132,N198,N396,N462,N67,N134,N201,N402,N469,N68,N136,N204,N408,N476,N69,N138,N207,N414,N483,N70,N140,N210,N420,N490,N71,N142,N213,N426,N497,N72,N144,N216,N432,N504,N73,N146,N219,N438,N511,N74,N148,N222,N444,N518,N75,N150,N225,N450,N525,N76,N152,N228,N456,N532,N77,N154,N231,N462,N539,N78,N156,N234,N468,N546,N79,N158,N237,N474,N553,N80,N160,N240,N480,N560,N81,N162,N243,N486,N567,N82,N164,N246,N492,N574,N83,N166,N249,N498,N581,N84,N168,N252,N504,N588,N85,N170,N255,N510,N595,N86,N172,N258,N516,N602,N87,N174,N261,N522,N609,N88,N176,N264,N528,N616,N89,N178,N267,N534,N623,N90,N180,N270,N540,N630,N91,N182,N273,N546,N637,N92,N184,N276,N552,N644,N93,N186,N279,N558,N651,N94,N188,N282,N564,N658,N95,N190,N285,N570,N665,N96,N192,N288,N576,N672,N97,N194,N291,N582,N679,N98,N196,N294,N588,N686,N99,N198,N297,N594,N693,N100,N200,N300,N600,N700,N101,N202,N303,N606,N707,N102,N204,N306,N612,N714,N103,N206,N309,N618,N721,N104,N208,N312,N624,N728,N105,N210,N315,N630,N735,N106,N212,N318,N636,N742,N107,N214,N321,N642,N749,N108,N216,N324,N648,N756,N109,N218,N327,N654,N763,N110,N220,N330,N660,N770,N111,N222,N333,N666,N777,N112,N224,N336,N672,N784,N113,N226,N339,N678,N791,N114,N228,N342,N684,N798,N115,N230,N345,N690,N805,N116,N232,N348,N696,N812,N117,N234,N351,N702,N819,N118,N236,N354,N708,N826,N119,N238,N357,N714,N833,N120,N240,N360,N720,N840,N121,N242,N363,N726,N847,N122,N244,N366,N732,N854,N123,N246,N369,N738,N861,N124,N248,N372,N744,N868,N125,N250,N375,N750,N875,N126,N252,N378,N756,N882,N127,N254,N381,N762,N889,N128,N256,N384,N768,N896,N129,N258,N387,N774,N903,N130,N260,N390,N780,N910,N131,N262,N393,N786,N917,N132,N264,N396,N792,N924,N133,N266,N399,N798,N931,N134,N268,N402,N804,N938,N135,N270,N405,N810,N945,N136,N272,N408,N816,N952,N137,N274,N411,N822,N959,N138,N276,N414,N828,N966,N139,N278,N417,N834,N973,N140,N280,N420,N840,N980,N141,N282,N423,N846,N987,N142,N284,N426,N852,N994,N143,N286,N429,N858,N1001,N144,N288,N432,N864,N1008,N145,N290,N435,N870,N1015,N146,N292,N438,N876,N1022,N147,N294,N441,N882,N1029,N148,N296,N444,N888,N1036,N149,N298,N447,N894,N1043,N150,N300,N450,N900,N1050,N151,N302,N453,N906,N1057,N152,N304,N456,N912,N1064,N153,N306,N459,N918,N1071,N154,N308,N462,N924,N1078,N155,N310,N465,N930,N1085,N156,N312,N468,N936,N1092,N157,N314,N471,N942,N1099,N158,N316,N474,N948,N1106,N159,N318,N477,N954,N1113,N160,N320,N480,N960,N1120,N161,N322,N483,N966,N1127,N162,N324,N486,N972,N1134,N163,N326,N489,N978,N1141,N164,N328,N492,N984,N1148,N165,N330,N495,N990,N1155,N166,N332,N498,N996,N1162,N167,N334,N501,N1002,N1169,N168,N336,N504,N1008,N1176,N169,N338,N507,N1014,N1183,N170,N340,N510,N1020,N1190,N171,N342,N513,N1026,N1197,N172,N344,N516,N1032,N1204,N173,N346,N519,N1038,N1211,N174,N348,N522,N1044,N1218,N175,N350,N525,N1050,N1225,N176,N352,N528,N1056,N1232,N177,N354,N531,N1062,N1239,N178,N356,N534,N1068,N1246,N179,N358,N537,N1074,N1253,N180,N360,N540,N1080,N1260,N181,N362,N543,N1086,N1267,N182,N364,N546,N1092,N1274,N183,N366,N549,N1098,N1281,N184,N368,N552,N1104,N1288,N185,N370,N555,N1110,N1295,N186,N372,N558,N1116,N1302,N187,N374,N561,N1122,N1309,N188,N376,N564,N1128,N1316,N189,N378,N567,N1134,N1323,N190,N380,N570,N1140,N1330,N191,N382,N573,N1146,N1337,N192,N384,N576,N1152,N1344,N193,N386,N579,N1158,N1351,N194,N388,N582,N1164,N1358,N195,N390,N585,N1170,N1365,N196,N392,N588,N1176,N1372,N197,N394,N591,N1182,N1379,N198,N396,N594,N1188,N1386,N199,N398,N597,N1194,N1393,N200,N400,N600,N1200,N1400,N201,N402,N603,N1206,N1407,N202,N404,N606,N1212,N1414,N203,N406,N609,N1218,N1421,N204,N408,N612,N1224,N1428,N205,N410,N615,N1230,N1435,N206,N412,N618,N1236,N1442,N207,N414,N621,N1242,N1449,N208,N416,N624,N1248,N1456,N209,N418,N627,N1254,N1463,N210,N420,N630,N1260,N1470,N211,N422,N633,N1266,N1477,N212,N424,N636,N1272,N1484,N213,N426,N639,N1278,N1491,N214,N428,N642,N1284,N1498,N215,N430,N645,N1290,N1505,N216,N432,N648,N1296,N1512,N217,N434,N651,N1302,N1519,N218,N436,N654,N1308,N1526,N219,N438,N657,N1314,N1533,N220,N440,N660,N1320,N1540,N221,N442,N663,N1326,N1547,N222,N444,N666,N1332,N1554,N223,N446,N669,N1338,N1561,N224,N448,N672,N1344,N1568,N225,N450,N675,N1350,N1575,N226,N452,N678,N1356,N1582,N227,N454,N681,N1362,N1589,N228,N456,N684,N1368,N1596,N229,N458,N687,N1374,N1603,N230,N460,N690,N1380,N1610,N231,N462,N693,N1386,N1617,N232,N464,N696,N1392,N1624,N233,N466,N699,N1398,N1631,N234,N468,N702,N1404,N1638,N235,N470,N705,N1410,N1645,N236,N472,N708,N1416,N1652,N237,N474,N711,N1422,N1659,N238,N476,N714,N1428,N1666,N239,N478,N717,N1434,N1673,N240,N480,N720,N1440,N1680,N241,N482,N723,N1446,N1687,N242,N484,N726,N1452,N1694,N243,N486,N729,N1458,N1701,N244,N488,N732,N1464,N1708,N245,N490,N735,N1470,N1715,N246,N492,N738,N1476,N1722,N247,N494,N741,N1482,N1729,N248,N496,N744,N1488,N1736,N249,N498,N747,N1494,N1743,N250,N500,N750,N1500,N1750,N251,N502,N753,N1506,N1757,N252,N504,N756,N1512,N1764,N253,N506,N759,N1518,N1771,N254,N508,N762,N1524,N1778,N255,N510,N765,N1530,N1785,N256,N512,N768,N1536,N1792,N257,N514,N771,N1542,N1799,N258,N516,N774,N1548,N1806,N259,N518,N777,N1554,N1813,N260,N520,N780,N1560,N1820,N261,N522,N783,N1566,N1827,N262,N524,N786,N1572,N1834,N263,N526,N789,N1578,N1841,N264,N528,N792,N1584,N1848,N265,N530,N795,N1590,N1855,N22,N23,N374,N391,N396,N414,N418,N437,N440,N460,N462,N483,N484,N506,N506,N529,N528,N552,N550,N575,N572,N598,N594,N621,N616,N644,N638,N667,N660,N690,N682,N713,N704,N736,N726,N759,N748,N782,N770,N805,N792,N828,N814,N851,N836,N874,N858,N897,N880,N920,N902,N943,N924,N966,N946,N989,N968,N1012,N990,N1035,N1012,N1058,N1034,N1081,N1056,N1104,N1078,N1127,N1100,N1150,N1122,N1173,N1144,N1196,N1166,N1219,N1188,N1242,N1210,N1265,N1232,N1288,N1254,N1311,N1276,N1334,N1298,N1357,N1320,N1380,N1342,N1403,N1364,N1426,N1386,N1449,N1408,N1472,N1430,N1495,N1452,N1518,N1474,N1541,N1496,N1564,N1518,N1587,N1540,N1610,N1562,N1633,N1584,N1656,N1606,N1679,N1628,N1702,N1650,N1725,N1672,N1748,N1694,N1771,N1716,N1794,N1738,N1817,N1760,N1840,N1782,N1863,N1804,N1886,N1826,N1909,N1848,N1932,N1870,N1955,N1892,N1978,N1914,N2001,N1936,N2024,N1958,N2047,N1980,N2070,N2002,N2093,N2024,N2116,N2046,N2139,N2068,N2162,N2090,N2185,N2112,N2208,N2134,N2231,N2156,N2254,N2178,N2277,N2200,N2300,N2222,N2323,N2244,N2346,N2266,N2369,N2288,N2392,N2310,N2415,N2332,N2438,N2354,N2461,N2376,N2484,N2398,N2507,N2420,N2530,N2442,N2553,N2464,N2576,N2486,N2599,N2508,N2622,N2530,N2645,N2552,N2668,N2574,N2691,N2596,N2714,N2618,N2737,N2640,N2760,N2662,N2783,N2684,N2806,N2706,N2829,N2728,N2852,N2750,N2875,N2772,N2898,N2794,N2921,N2816,N2944,N2838,N2967,N2860,N2990,N2882,N3013,N2904,N3036,N2926,N3059,N2948,N3082,N2970,N3105,N2992,N3128,N3014,N3151,N3036,N3174,N3058,N3197,N3080,N3220,N3102,N3243,N3124,N3266,N3146,N3289,N3168,N3312,N3190,N3335,N3212,N3358,N3234,N3381,N3256,N3404,N3278,N3427,N3300,N3450,N3322,N3473,N3344,N3496,N3366,N3519,N3388,N3542,N3410,N3565,N3432,N3588,N3454,N3611,N3476,N3634,N3498,N3657,N3520,N3680,N3542,N3703,N3564,N3726,N3586,N3749,N3608,N3772,N3630,N3795,N3652,N3818,N3674,N3841,N3696,N3864,N3718,N3887,N3740,N3910,N3762,N3933,N3784,N3956,N3806,N3979,N3828,N4002,N3850,N4025,N3872,N4048,N3894,N4071,N3916,N4094,N3938,N4117,N3960,N4140,N3982,N4163,N4004,N4186,N4026,N4209,N4048,N4232,N4070,N4255,N4092,N4278,N4114,N4301,N4136,N4324,N4158,N4347,N4180,N4370,N4202,N4393,N4224,N4416,N4246,N4439,N4268,N4462,N4290,N4485,N4312,N4508,N4334,N4531,N4356,N4554,N4378,N4577,N4400,N4600,N4422,N4623,N4444,N4646,N4466,N4669,N4488,N4692,N4510,N4715,N4532,N4738,N4554,N4761,N4576,N4784,N4598,N4807,N4620,N4830,N4642,N4853,N4664,N4876,N4686,N4899,N4708,N4922,N4730,N4945,N4752,N4968,N4774,N4991,N4796,N5014,N4818,N5037,N4840,N5060,N4862,N5083,N4884,N5106,N4906,N5129,N4928,N5152,N4950,N5175,N4972,N5198,N4994,N5221,N5016,N5244,N5038,N5267,N5060,N5290,N5082,N5313,N5104,N5336,N5126,N5359,N5148,N5382,N5170,N5405,N5192,N5428,N5214,N5451,N5236,N5474,N5258,N5497,N5280,N5520,N5302,N5543,N5324,N5566,N5346,N5589,N5368,N5612,N5390,N5635,N5412,N5658,N5434,N5681,N5456,N5704,N5478,N5727,N5500,N5750,N5522,N5773,N5544,N5796,N5566,N5819,N5588,N5842,N5610,N5865,N5632,N5888,N5654,N5911,N5676,N5934,N5698,N5957,N5720,N5980,N5742,N6003,N5764,N6026,N5786,N6049,N5808,N6072,N5830,N6095);

input N1,N2,N3,N6,N7,N17,N34,N51,N102,N119,N18,N36,N54,N108,N126,N19,N38,N57,N114,N133,N20,N40,N60,N120,N140,N21,N42,N63,N126,N147,N22,N44,N66,N132,N154,N23,N46,N69,N138,N161,N24,N48,N72,N144,N168,N25,N50,N75,N150,N175,N26,N52,N78,N156,N182,N27,N54,N81,N162,N189,N28,N56,N84,N168,N196,N29,N58,N87,N174,N203,N30,N60,N90,N180,N210,N31,N62,N93,N186,N217,N32,N64,N96,N192,N224,N33,N66,N99,N198,N231,N34,N68,N102,N204,N238,N35,N70,N105,N210,N245,N36,N72,N108,N216,N252,N37,N74,N111,N222,N259,N38,N76,N114,N228,N266,N39,N78,N117,N234,N273,N40,N80,N120,N240,N280,N41,N82,N123,N246,N287,N42,N84,N126,N252,N294,N43,N86,N129,N258,N301,N44,N88,N132,N264,N308,N45,N90,N135,N270,N315,N46,N92,N138,N276,N322,N47,N94,N141,N282,N329,N48,N96,N144,N288,N336,N49,N98,N147,N294,N343,N50,N100,N150,N300,N350,N51,N102,N153,N306,N357,N52,N104,N156,N312,N364,N53,N106,N159,N318,N371,N54,N108,N162,N324,N378,N55,N110,N165,N330,N385,N56,N112,N168,N336,N392,N57,N114,N171,N342,N399,N58,N116,N174,N348,N406,N59,N118,N177,N354,N413,N60,N120,N180,N360,N420,N61,N122,N183,N366,N427,N62,N124,N186,N372,N434,N63,N126,N189,N378,N441,N64,N128,N192,N384,N448,N65,N130,N195,N390,N455,N66,N132,N198,N396,N462,N67,N134,N201,N402,N469,N68,N136,N204,N408,N476,N69,N138,N207,N414,N483,N70,N140,N210,N420,N490,N71,N142,N213,N426,N497,N72,N144,N216,N432,N504,N73,N146,N219,N438,N511,N74,N148,N222,N444,N518,N75,N150,N225,N450,N525,N76,N152,N228,N456,N532,N77,N154,N231,N462,N539,N78,N156,N234,N468,N546,N79,N158,N237,N474,N553,N80,N160,N240,N480,N560,N81,N162,N243,N486,N567,N82,N164,N246,N492,N574,N83,N166,N249,N498,N581,N84,N168,N252,N504,N588,N85,N170,N255,N510,N595,N86,N172,N258,N516,N602,N87,N174,N261,N522,N609,N88,N176,N264,N528,N616,N89,N178,N267,N534,N623,N90,N180,N270,N540,N630,N91,N182,N273,N546,N637,N92,N184,N276,N552,N644,N93,N186,N279,N558,N651,N94,N188,N282,N564,N658,N95,N190,N285,N570,N665,N96,N192,N288,N576,N672,N97,N194,N291,N582,N679,N98,N196,N294,N588,N686,N99,N198,N297,N594,N693,N100,N200,N300,N600,N700,N101,N202,N303,N606,N707,N102,N204,N306,N612,N714,N103,N206,N309,N618,N721,N104,N208,N312,N624,N728,N105,N210,N315,N630,N735,N106,N212,N318,N636,N742,N107,N214,N321,N642,N749,N108,N216,N324,N648,N756,N109,N218,N327,N654,N763,N110,N220,N330,N660,N770,N111,N222,N333,N666,N777,N112,N224,N336,N672,N784,N113,N226,N339,N678,N791,N114,N228,N342,N684,N798,N115,N230,N345,N690,N805,N116,N232,N348,N696,N812,N117,N234,N351,N702,N819,N118,N236,N354,N708,N826,N119,N238,N357,N714,N833,N120,N240,N360,N720,N840,N121,N242,N363,N726,N847,N122,N244,N366,N732,N854,N123,N246,N369,N738,N861,N124,N248,N372,N744,N868,N125,N250,N375,N750,N875,N126,N252,N378,N756,N882,N127,N254,N381,N762,N889,N128,N256,N384,N768,N896,N129,N258,N387,N774,N903,N130,N260,N390,N780,N910,N131,N262,N393,N786,N917,N132,N264,N396,N792,N924,N133,N266,N399,N798,N931,N134,N268,N402,N804,N938,N135,N270,N405,N810,N945,N136,N272,N408,N816,N952,N137,N274,N411,N822,N959,N138,N276,N414,N828,N966,N139,N278,N417,N834,N973,N140,N280,N420,N840,N980,N141,N282,N423,N846,N987,N142,N284,N426,N852,N994,N143,N286,N429,N858,N1001,N144,N288,N432,N864,N1008,N145,N290,N435,N870,N1015,N146,N292,N438,N876,N1022,N147,N294,N441,N882,N1029,N148,N296,N444,N888,N1036,N149,N298,N447,N894,N1043,N150,N300,N450,N900,N1050,N151,N302,N453,N906,N1057,N152,N304,N456,N912,N1064,N153,N306,N459,N918,N1071,N154,N308,N462,N924,N1078,N155,N310,N465,N930,N1085,N156,N312,N468,N936,N1092,N157,N314,N471,N942,N1099,N158,N316,N474,N948,N1106,N159,N318,N477,N954,N1113,N160,N320,N480,N960,N1120,N161,N322,N483,N966,N1127,N162,N324,N486,N972,N1134,N163,N326,N489,N978,N1141,N164,N328,N492,N984,N1148,N165,N330,N495,N990,N1155,N166,N332,N498,N996,N1162,N167,N334,N501,N1002,N1169,N168,N336,N504,N1008,N1176,N169,N338,N507,N1014,N1183,N170,N340,N510,N1020,N1190,N171,N342,N513,N1026,N1197,N172,N344,N516,N1032,N1204,N173,N346,N519,N1038,N1211,N174,N348,N522,N1044,N1218,N175,N350,N525,N1050,N1225,N176,N352,N528,N1056,N1232,N177,N354,N531,N1062,N1239,N178,N356,N534,N1068,N1246,N179,N358,N537,N1074,N1253,N180,N360,N540,N1080,N1260,N181,N362,N543,N1086,N1267,N182,N364,N546,N1092,N1274,N183,N366,N549,N1098,N1281,N184,N368,N552,N1104,N1288,N185,N370,N555,N1110,N1295,N186,N372,N558,N1116,N1302,N187,N374,N561,N1122,N1309,N188,N376,N564,N1128,N1316,N189,N378,N567,N1134,N1323,N190,N380,N570,N1140,N1330,N191,N382,N573,N1146,N1337,N192,N384,N576,N1152,N1344,N193,N386,N579,N1158,N1351,N194,N388,N582,N1164,N1358,N195,N390,N585,N1170,N1365,N196,N392,N588,N1176,N1372,N197,N394,N591,N1182,N1379,N198,N396,N594,N1188,N1386,N199,N398,N597,N1194,N1393,N200,N400,N600,N1200,N1400,N201,N402,N603,N1206,N1407,N202,N404,N606,N1212,N1414,N203,N406,N609,N1218,N1421,N204,N408,N612,N1224,N1428,N205,N410,N615,N1230,N1435,N206,N412,N618,N1236,N1442,N207,N414,N621,N1242,N1449,N208,N416,N624,N1248,N1456,N209,N418,N627,N1254,N1463,N210,N420,N630,N1260,N1470,N211,N422,N633,N1266,N1477,N212,N424,N636,N1272,N1484,N213,N426,N639,N1278,N1491,N214,N428,N642,N1284,N1498,N215,N430,N645,N1290,N1505,N216,N432,N648,N1296,N1512,N217,N434,N651,N1302,N1519,N218,N436,N654,N1308,N1526,N219,N438,N657,N1314,N1533,N220,N440,N660,N1320,N1540,N221,N442,N663,N1326,N1547,N222,N444,N666,N1332,N1554,N223,N446,N669,N1338,N1561,N224,N448,N672,N1344,N1568,N225,N450,N675,N1350,N1575,N226,N452,N678,N1356,N1582,N227,N454,N681,N1362,N1589,N228,N456,N684,N1368,N1596,N229,N458,N687,N1374,N1603,N230,N460,N690,N1380,N1610,N231,N462,N693,N1386,N1617,N232,N464,N696,N1392,N1624,N233,N466,N699,N1398,N1631,N234,N468,N702,N1404,N1638,N235,N470,N705,N1410,N1645,N236,N472,N708,N1416,N1652,N237,N474,N711,N1422,N1659,N238,N476,N714,N1428,N1666,N239,N478,N717,N1434,N1673,N240,N480,N720,N1440,N1680,N241,N482,N723,N1446,N1687,N242,N484,N726,N1452,N1694,N243,N486,N729,N1458,N1701,N244,N488,N732,N1464,N1708,N245,N490,N735,N1470,N1715,N246,N492,N738,N1476,N1722,N247,N494,N741,N1482,N1729,N248,N496,N744,N1488,N1736,N249,N498,N747,N1494,N1743,N250,N500,N750,N1500,N1750,N251,N502,N753,N1506,N1757,N252,N504,N756,N1512,N1764,N253,N506,N759,N1518,N1771,N254,N508,N762,N1524,N1778,N255,N510,N765,N1530,N1785,N256,N512,N768,N1536,N1792,N257,N514,N771,N1542,N1799,N258,N516,N774,N1548,N1806,N259,N518,N777,N1554,N1813,N260,N520,N780,N1560,N1820,N261,N522,N783,N1566,N1827,N262,N524,N786,N1572,N1834,N263,N526,N789,N1578,N1841,N264,N528,N792,N1584,N1848,N265,N530,N795,N1590,N1855;

output N22,N23,N374,N391,N396,N414,N418,N437,N440,N460,N462,N483,N484,N506,N506,N529,N528,N552,N550,N575,N572,N598,N594,N621,N616,N644,N638,N667,N660,N690,N682,N713,N704,N736,N726,N759,N748,N782,N770,N805,N792,N828,N814,N851,N836,N874,N858,N897,N880,N920,N902,N943,N924,N966,N946,N989,N968,N1012,N990,N1035,N1012,N1058,N1034,N1081,N1056,N1104,N1078,N1127,N1100,N1150,N1122,N1173,N1144,N1196,N1166,N1219,N1188,N1242,N1210,N1265,N1232,N1288,N1254,N1311,N1276,N1334,N1298,N1357,N1320,N1380,N1342,N1403,N1364,N1426,N1386,N1449,N1408,N1472,N1430,N1495,N1452,N1518,N1474,N1541,N1496,N1564,N1518,N1587,N1540,N1610,N1562,N1633,N1584,N1656,N1606,N1679,N1628,N1702,N1650,N1725,N1672,N1748,N1694,N1771,N1716,N1794,N1738,N1817,N1760,N1840,N1782,N1863,N1804,N1886,N1826,N1909,N1848,N1932,N1870,N1955,N1892,N1978,N1914,N2001,N1936,N2024,N1958,N2047,N1980,N2070,N2002,N2093,N2024,N2116,N2046,N2139,N2068,N2162,N2090,N2185,N2112,N2208,N2134,N2231,N2156,N2254,N2178,N2277,N2200,N2300,N2222,N2323,N2244,N2346,N2266,N2369,N2288,N2392,N2310,N2415,N2332,N2438,N2354,N2461,N2376,N2484,N2398,N2507,N2420,N2530,N2442,N2553,N2464,N2576,N2486,N2599,N2508,N2622,N2530,N2645,N2552,N2668,N2574,N2691,N2596,N2714,N2618,N2737,N2640,N2760,N2662,N2783,N2684,N2806,N2706,N2829,N2728,N2852,N2750,N2875,N2772,N2898,N2794,N2921,N2816,N2944,N2838,N2967,N2860,N2990,N2882,N3013,N2904,N3036,N2926,N3059,N2948,N3082,N2970,N3105,N2992,N3128,N3014,N3151,N3036,N3174,N3058,N3197,N3080,N3220,N3102,N3243,N3124,N3266,N3146,N3289,N3168,N3312,N3190,N3335,N3212,N3358,N3234,N3381,N3256,N3404,N3278,N3427,N3300,N3450,N3322,N3473,N3344,N3496,N3366,N3519,N3388,N3542,N3410,N3565,N3432,N3588,N3454,N3611,N3476,N3634,N3498,N3657,N3520,N3680,N3542,N3703,N3564,N3726,N3586,N3749,N3608,N3772,N3630,N3795,N3652,N3818,N3674,N3841,N3696,N3864,N3718,N3887,N3740,N3910,N3762,N3933,N3784,N3956,N3806,N3979,N3828,N4002,N3850,N4025,N3872,N4048,N3894,N4071,N3916,N4094,N3938,N4117,N3960,N4140,N3982,N4163,N4004,N4186,N4026,N4209,N4048,N4232,N4070,N4255,N4092,N4278,N4114,N4301,N4136,N4324,N4158,N4347,N4180,N4370,N4202,N4393,N4224,N4416,N4246,N4439,N4268,N4462,N4290,N4485,N4312,N4508,N4334,N4531,N4356,N4554,N4378,N4577,N4400,N4600,N4422,N4623,N4444,N4646,N4466,N4669,N4488,N4692,N4510,N4715,N4532,N4738,N4554,N4761,N4576,N4784,N4598,N4807,N4620,N4830,N4642,N4853,N4664,N4876,N4686,N4899,N4708,N4922,N4730,N4945,N4752,N4968,N4774,N4991,N4796,N5014,N4818,N5037,N4840,N5060,N4862,N5083,N4884,N5106,N4906,N5129,N4928,N5152,N4950,N5175,N4972,N5198,N4994,N5221,N5016,N5244,N5038,N5267,N5060,N5290,N5082,N5313,N5104,N5336,N5126,N5359,N5148,N5382,N5170,N5405,N5192,N5428,N5214,N5451,N5236,N5474,N5258,N5497,N5280,N5520,N5302,N5543,N5324,N5566,N5346,N5589,N5368,N5612,N5390,N5635,N5412,N5658,N5434,N5681,N5456,N5704,N5478,N5727,N5500,N5750,N5522,N5773,N5544,N5796,N5566,N5819,N5588,N5842,N5610,N5865,N5632,N5888,N5654,N5911,N5676,N5934,N5698,N5957,N5720,N5980,N5742,N6003,N5764,N6026,N5786,N6049,N5808,N6072,N5830,N6095;

wire N10,N11,N16,N19,N170,N187,N272,N323,N180,N198,N288,N342,N190,N209,N304,N361,N200,N220,N320,N380,N210,N231,N336,N399,N220,N242,N352,N230,N253,N368,N240,N264,N384,N456,N250,N275,N400,N475,N260,N286,N416,N494,N270,N297,N432,N513,N280,N308,N448,N532,N290,N319,N464,N551,N300,N330,N480,N570,N310,N341,N496,N589,N320,N352,N512,N608,N330,N363,N627,N340,N544,N646,N350,N385,N560,N665,N360,N576,N684,N370,N407,N592,N703,N380,N608,N722,N390,N429,N624,N741,N400,N640,N760,N410,N451,N656,N779,N420,N672,N798,N430,N473,N688,N817,N450,N495,N720,N855,N470,N517,N752,N893,N480,N768,N912,N490,N539,N784,N931,N500,N800,N950,N510,N561,N816,N969,N520,N832,N988,N530,N583,N848,N1007,N540,N864,N1026,N605,N1045,N560,N896,N1064,N570,N627,N912,N1083,N580,N928,N1102,N590,N649,N944,N1121,N600,N960,N1140,N610,N671,N976,N1159,N620,N992,N1178,N630,N693,N1008,N1197,N640,N1024,N1216,N650,N715,N1040,N1235,N670,N737,N1072,N1273,N680,N1088,N1292,N700,N1120,N1330,N710,N781,N1136,N1349,N720,N1152,N1368,N730,N803,N1168,N1387,N740,N1184,N1406,N750,N825,N1200,N1425,N760,N1216,N1444,N847,N1463,N780,N1248,N1482,N790,N869,N1264,N1501,N800,N1280,N1520,N810,N891,N1296,N1539,N820,N1312,N1558,N830,N913,N1328,N1577,N840,N1344,N1596,N850,N935,N1360,N1615,N860,N1376,N1634,N870,N957,N1392,N1653,N890,N979,N1424,N1691,N900,N1440,N1710,N910,N1001,N1456,N1729,N930,N1023,N1488,N1767,N940,N1504,N1786,N950,N1045,N1520,N1805,N960,N1536,N1824,N970,N1067,N1552,N1843,N980,N1568,N1862,N1089,N1881,N1000,N1600,N1900,N1010,N1111,N1616,N1919,N1020,N1632,N1938,N1030,N1133,N1648,N1957,N1040,N1664,N1976,N1050,N1155,N1680,N1995,N1060,N1696,N2014,N1070,N1177,N1712,N2033,N1080,N1728,N2052,N1090,N1199,N1744,N2071,N1110,N1221,N1776,N2109,N1120,N1792,N2128,N1130,N1243,N1808,N2147,N1140,N1824,N2166,N1160,N1856,N2204,N1170,N1287,N1872,N2223,N1180,N1888,N2242,N1190,N1309,N1904,N2261,N1200,N1920,N2280,N1331,N2299,N1220,N1952,N2318,N1230,N1353,N1968,N2337,N1240,N1984,N2356,N1250,N1375,N2000,N2375,N1260,N2016,N2394,N1270,N1397,N2032,N2413,N1280,N2048,N2432,N1290,N1419,N2064,N2451,N1300,N2080,N2470,N1310,N1441,N2096,N2489,N1330,N1463,N2128,N2527,N1340,N2144,N2546,N1350,N1485,N2160,N2565,N1360,N2176,N2584,N1370,N1507,N2192,N2603,N1390,N1529,N2224,N2641,N1400,N2240,N2660,N1410,N1551,N2256,N2679,N1420,N2272,N2698,N1573,N2717,N1440,N2304,N2736,N1450,N1595,N2320,N2755,N1460,N2336,N2774,N1470,N1617,N2352,N2793,N1480,N2368,N2812,N1490,N1639,N2384,N2831,N1500,N2400,N2850,N1510,N1661,N2416,N2869,N1520,N2432,N2888,N1530,N1683,N2448,N2907,N1550,N1705,N2480,N2945,N1560,N2496,N2964,N1570,N1727,N2512,N2983,N1580,N2528,N3002,N1590,N1749,N2544,N3021,N1600,N2560,N3040,N1620,N2592,N3078,N1630,N1793,N2608,N3097,N1640,N2624,N3116,N1815,N3135,N1660,N2656,N3154,N1670,N1837,N2672,N3173,N1680,N2688,N3192,N1690,N1859,N2704,N3211,N1700,N2720,N3230,N1710,N1881,N2736,N3249,N1720,N2752,N3268,N1730,N1903,N2768,N3287,N1740,N2784,N3306,N1750,N1925,N2800,N3325,N1770,N1947,N2832,N3363,N1780,N2848,N3382,N1790,N1969,N2864,N3401,N1800,N2880,N3420,N1810,N1991,N2896,N3439,N1820,N2912,N3458;

nand NAND2_1 (N10, N1616, N4092);
nand NAND2_2 (N11, N1919, N4278);
nand NAND2_3 (N16, N2222, N1870);
nand NAND2_4 (N19, N2323, N2057);
nand NAND2_5 (N22, N1020, N2992);
nand NAND2_6 (N23, N1122, N3553);
nand NAND2_7 (N170, N1632, N4114);
nand NAND2_8 (N187, N1938, N4301);
nand NAND2_9 (N272, N2244, N1880);
nand NAND2_10 (N323, N2346, N2068);
nand NAND2_11 (N374, N1030, N3008);
nand NAND2_12 (N391, N1133, N3572);
nand NAND2_13 (N180, N1648, N4136);
nand NAND2_14 (N198, N1957, N4324);
nand NAND2_15 (N288, N2266, N1890);
nand NAND2_16 (N342, N2369, N2079);
nand NAND2_17 (N396, N1040, N3024);
nand NAND2_18 (N414, N1144, N3591);
nand NAND2_19 (N190, N1664, N4158);
nand NAND2_20 (N209, N1976, N4347);
nand NAND2_21 (N304, N2288, N1900);
nand NAND2_22 (N361, N2392, N2090);
nand NAND2_23 (N418, N1050, N3040);
nand NAND2_24 (N437, N1155, N3610);
nand NAND2_25 (N200, N1680, N4180);
nand NAND2_26 (N220, N1995, N4370);
nand NAND2_27 (N320, N2310, N1910);
nand NAND2_28 (N380, N2415, N2101);
nand NAND2_29 (N440, N1060, N3056);
nand NAND2_30 (N460, N1166, N3629);
nand NAND2_31 (N210, N1696, N4202);
nand NAND2_32 (N231, N2014, N4393);
nand NAND2_33 (N336, N2332, N1920);
nand NAND2_34 (N399, N2438, N2112);
nand NAND2_35 (N462, N1070, N3072);
nand NAND2_36 (N483, N1177, N3648);
nand NAND2_37 (N220, N1712, N4224);
nand NAND2_38 (N242, N2033, N4416);
nand NAND2_39 (N352, N2354, N1930);
nand NAND2_40 (N418, N2461, N2123);
nand NAND2_41 (N484, N1080, N3088);
nand NAND2_42 (N506, N1188, N3667);
nand NAND2_43 (N230, N1728, N4246);
nand NAND2_44 (N253, N2052, N4439);
nand NAND2_45 (N368, N2376, N1940);
nand NAND2_46 (N437, N2484, N2134);
nand NAND2_47 (N506, N1090, N3104);
nand NAND2_48 (N529, N1199, N3686);
nand NAND2_49 (N240, N1744, N4268);
nand NAND2_50 (N264, N2071, N4462);
nand NAND2_51 (N384, N2398, N1950);
nand NAND2_52 (N456, N2507, N2145);
nand NAND2_53 (N528, N1100, N3120);
nand NAND2_54 (N552, N1210, N3705);
nand NAND2_55 (N250, N1760, N4290);
nand NAND2_56 (N275, N2090, N4485);
nand NAND2_57 (N400, N2420, N1960);
nand NAND2_58 (N475, N2530, N2156);
nand NAND2_59 (N550, N1110, N3136);
nand NAND2_60 (N575, N1221, N3724);
nand NAND2_61 (N260, N1776, N4312);
nand NAND2_62 (N286, N2109, N4508);
nand NAND2_63 (N416, N2442, N1970);
nand NAND2_64 (N494, N2553, N2167);
nand NAND2_65 (N572, N1120, N3152);
nand NAND2_66 (N598, N1232, N3743);
nand NAND2_67 (N270, N1792, N4334);
nand NAND2_68 (N297, N2128, N4531);
nand NAND2_69 (N432, N2464, N1980);
nand NAND2_70 (N513, N2576, N2178);
nand NAND2_71 (N594, N1130, N3168);
nand NAND2_72 (N621, N1243, N3762);
nand NAND2_73 (N280, N1808, N4356);
nand NAND2_74 (N308, N2147, N4554);
nand NAND2_75 (N448, N2486, N1990);
nand NAND2_76 (N532, N2599, N2189);
nand NAND2_77 (N616, N1140, N3184);
nand NAND2_78 (N644, N1254, N3781);
nand NAND2_79 (N290, N1824, N4378);
nand NAND2_80 (N319, N2166, N4577);
nand NAND2_81 (N464, N2508, N2000);
nand NAND2_82 (N551, N2622, N2200);
nand NAND2_83 (N638, N1150, N3200);
nand NAND2_84 (N667, N1265, N3800);
nand NAND2_85 (N300, N1840, N4400);
nand NAND2_86 (N330, N2185, N4600);
nand NAND2_87 (N480, N2530, N2010);
nand NAND2_88 (N570, N2645, N2211);
nand NAND2_89 (N660, N1160, N3216);
nand NAND2_90 (N690, N1276, N3819);
nand NAND2_91 (N310, N1856, N4422);
nand NAND2_92 (N341, N2204, N4623);
nand NAND2_93 (N496, N2552, N2020);
nand NAND2_94 (N589, N2668, N2222);
nand NAND2_95 (N682, N1170, N3232);
nand NAND2_96 (N713, N1287, N3838);
nand NAND2_97 (N320, N1872, N4444);
nand NAND2_98 (N352, N2223, N4646);
nand NAND2_99 (N512, N2574, N2030);
nand NAND2_100 (N608, N2691, N2233);
nand NAND2_101 (N704, N1180, N3248);
nand NAND2_102 (N736, N1298, N3857);
nand NAND2_103 (N330, N1888, N4466);
nand NAND2_104 (N363, N2242, N4669);
nand NAND2_105 (N528, N2596, N2040);
nand NAND2_106 (N627, N2714, N2244);
nand NAND2_107 (N726, N1190, N3264);
nand NAND2_108 (N759, N1309, N3876);
nand NAND2_109 (N340, N1904, N4488);
nand NAND2_110 (N374, N2261, N4692);
nand NAND2_111 (N544, N2618, N2050);
nand NAND2_112 (N646, N2737, N2255);
nand NAND2_113 (N748, N1200, N3280);
nand NAND2_114 (N782, N1320, N3895);
nand NAND2_115 (N350, N1920, N4510);
nand NAND2_116 (N385, N2280, N4715);
nand NAND2_117 (N560, N2640, N2060);
nand NAND2_118 (N665, N2760, N2266);
nand NAND2_119 (N770, N1210, N3296);
nand NAND2_120 (N805, N1331, N3914);
nand NAND2_121 (N360, N1936, N4532);
nand NAND2_122 (N396, N2299, N4738);
nand NAND2_123 (N576, N2662, N2070);
nand NAND2_124 (N684, N2783, N2277);
nand NAND2_125 (N792, N1220, N3312);
nand NAND2_126 (N828, N1342, N3933);
nand NAND2_127 (N370, N1952, N4554);
nand NAND2_128 (N407, N2318, N4761);
nand NAND2_129 (N592, N2684, N2080);
nand NAND2_130 (N703, N2806, N2288);
nand NAND2_131 (N814, N1230, N3328);
nand NAND2_132 (N851, N1353, N3952);
nand NAND2_133 (N380, N1968, N4576);
nand NAND2_134 (N418, N2337, N4784);
nand NAND2_135 (N608, N2706, N2090);
nand NAND2_136 (N722, N2829, N2299);
nand NAND2_137 (N836, N1240, N3344);
nand NAND2_138 (N874, N1364, N3971);
nand NAND2_139 (N390, N1984, N4598);
nand NAND2_140 (N429, N2356, N4807);
nand NAND2_141 (N624, N2728, N2100);
nand NAND2_142 (N741, N2852, N2310);
nand NAND2_143 (N858, N1250, N3360);
nand NAND2_144 (N897, N1375, N3990);
nand NAND2_145 (N400, N2000, N4620);
nand NAND2_146 (N440, N2375, N4830);
nand NAND2_147 (N640, N2750, N2110);
nand NAND2_148 (N760, N2875, N2321);
nand NAND2_149 (N880, N1260, N3376);
nand NAND2_150 (N920, N1386, N4009);
nand NAND2_151 (N410, N2016, N4642);
nand NAND2_152 (N451, N2394, N4853);
nand NAND2_153 (N656, N2772, N2120);
nand NAND2_154 (N779, N2898, N2332);
nand NAND2_155 (N902, N1270, N3392);
nand NAND2_156 (N943, N1397, N4028);
nand NAND2_157 (N420, N2032, N4664);
nand NAND2_158 (N462, N2413, N4876);
nand NAND2_159 (N672, N2794, N2130);
nand NAND2_160 (N798, N2921, N2343);
nand NAND2_161 (N924, N1280, N3408);
nand NAND2_162 (N966, N1408, N4047);
nand NAND2_163 (N430, N2048, N4686);
nand NAND2_164 (N473, N2432, N4899);
nand NAND2_165 (N688, N2816, N2140);
nand NAND2_166 (N817, N2944, N2354);
nand NAND2_167 (N946, N1290, N3424);
nand NAND2_168 (N989, N1419, N4066);
nand NAND2_169 (N440, N2064, N4708);
nand NAND2_170 (N484, N2451, N4922);
nand NAND2_171 (N704, N2838, N2150);
nand NAND2_172 (N836, N2967, N2365);
nand NAND2_173 (N968, N1300, N3440);
nand NAND2_174 (N1012, N1430, N4085);
nand NAND2_175 (N450, N2080, N4730);
nand NAND2_176 (N495, N2470, N4945);
nand NAND2_177 (N720, N2860, N2160);
nand NAND2_178 (N855, N2990, N2376);
nand NAND2_179 (N990, N1310, N3456);
nand NAND2_180 (N1035, N1441, N4104);
nand NAND2_181 (N460, N2096, N4752);
nand NAND2_182 (N506, N2489, N4968);
nand NAND2_183 (N736, N2882, N2170);
nand NAND2_184 (N874, N3013, N2387);
nand NAND2_185 (N1012, N1320, N3472);
nand NAND2_186 (N1058, N1452, N4123);
nand NAND2_187 (N470, N2112, N4774);
nand NAND2_188 (N517, N2508, N4991);
nand NAND2_189 (N752, N2904, N2180);
nand NAND2_190 (N893, N3036, N2398);
nand NAND2_191 (N1034, N1330, N3488);
nand NAND2_192 (N1081, N1463, N4142);
nand NAND2_193 (N480, N2128, N4796);
nand NAND2_194 (N528, N2527, N5014);
nand NAND2_195 (N768, N2926, N2190);
nand NAND2_196 (N912, N3059, N2409);
nand NAND2_197 (N1056, N1340, N3504);
nand NAND2_198 (N1104, N1474, N4161);
nand NAND2_199 (N490, N2144, N4818);
nand NAND2_200 (N539, N2546, N5037);
nand NAND2_201 (N784, N2948, N2200);
nand NAND2_202 (N931, N3082, N2420);
nand NAND2_203 (N1078, N1350, N3520);
nand NAND2_204 (N1127, N1485, N4180);
nand NAND2_205 (N500, N2160, N4840);
nand NAND2_206 (N550, N2565, N5060);
nand NAND2_207 (N800, N2970, N2210);
nand NAND2_208 (N950, N3105, N2431);
nand NAND2_209 (N1100, N1360, N3536);
nand NAND2_210 (N1150, N1496, N4199);
nand NAND2_211 (N510, N2176, N4862);
nand NAND2_212 (N561, N2584, N5083);
nand NAND2_213 (N816, N2992, N2220);
nand NAND2_214 (N969, N3128, N2442);
nand NAND2_215 (N1122, N1370, N3552);
nand NAND2_216 (N1173, N1507, N4218);
nand NAND2_217 (N520, N2192, N4884);
nand NAND2_218 (N572, N2603, N5106);
nand NAND2_219 (N832, N3014, N2230);
nand NAND2_220 (N988, N3151, N2453);
nand NAND2_221 (N1144, N1380, N3568);
nand NAND2_222 (N1196, N1518, N4237);
nand NAND2_223 (N530, N2208, N4906);
nand NAND2_224 (N583, N2622, N5129);
nand NAND2_225 (N848, N3036, N2240);
nand NAND2_226 (N1007, N3174, N2464);
nand NAND2_227 (N1166, N1390, N3584);
nand NAND2_228 (N1219, N1529, N4256);
nand NAND2_229 (N540, N2224, N4928);
nand NAND2_230 (N594, N2641, N5152);
nand NAND2_231 (N864, N3058, N2250);
nand NAND2_232 (N1026, N3197, N2475);
nand NAND2_233 (N1188, N1400, N3600);
nand NAND2_234 (N1242, N1540, N4275);
nand NAND2_235 (N550, N2240, N4950);
nand NAND2_236 (N605, N2660, N5175);
nand NAND2_237 (N880, N3080, N2260);
nand NAND2_238 (N1045, N3220, N2486);
nand NAND2_239 (N1210, N1410, N3616);
nand NAND2_240 (N1265, N1551, N4294);
nand NAND2_241 (N560, N2256, N4972);
nand NAND2_242 (N616, N2679, N5198);
nand NAND2_243 (N896, N3102, N2270);
nand NAND2_244 (N1064, N3243, N2497);
nand NAND2_245 (N1232, N1420, N3632);
nand NAND2_246 (N1288, N1562, N4313);
nand NAND2_247 (N570, N2272, N4994);
nand NAND2_248 (N627, N2698, N5221);
nand NAND2_249 (N912, N3124, N2280);
nand NAND2_250 (N1083, N3266, N2508);
nand NAND2_251 (N1254, N1430, N3648);
nand NAND2_252 (N1311, N1573, N4332);
nand NAND2_253 (N580, N2288, N5016);
nand NAND2_254 (N638, N2717, N5244);
nand NAND2_255 (N928, N3146, N2290);
nand NAND2_256 (N1102, N3289, N2519);
nand NAND2_257 (N1276, N1440, N3664);
nand NAND2_258 (N1334, N1584, N4351);
nand NAND2_259 (N590, N2304, N5038);
nand NAND2_260 (N649, N2736, N5267);
nand NAND2_261 (N944, N3168, N2300);
nand NAND2_262 (N1121, N3312, N2530);
nand NAND2_263 (N1298, N1450, N3680);
nand NAND2_264 (N1357, N1595, N4370);
nand NAND2_265 (N600, N2320, N5060);
nand NAND2_266 (N660, N2755, N5290);
nand NAND2_267 (N960, N3190, N2310);
nand NAND2_268 (N1140, N3335, N2541);
nand NAND2_269 (N1320, N1460, N3696);
nand NAND2_270 (N1380, N1606, N4389);
nand NAND2_271 (N610, N2336, N5082);
nand NAND2_272 (N671, N2774, N5313);
nand NAND2_273 (N976, N3212, N2320);
nand NAND2_274 (N1159, N3358, N2552);
nand NAND2_275 (N1342, N1470, N3712);
nand NAND2_276 (N1403, N1617, N4408);
nand NAND2_277 (N620, N2352, N5104);
nand NAND2_278 (N682, N2793, N5336);
nand NAND2_279 (N992, N3234, N2330);
nand NAND2_280 (N1178, N3381, N2563);
nand NAND2_281 (N1364, N1480, N3728);
nand NAND2_282 (N1426, N1628, N4427);
nand NAND2_283 (N630, N2368, N5126);
nand NAND2_284 (N693, N2812, N5359);
nand NAND2_285 (N1008, N3256, N2340);
nand NAND2_286 (N1197, N3404, N2574);
nand NAND2_287 (N1386, N1490, N3744);
nand NAND2_288 (N1449, N1639, N4446);
nand NAND2_289 (N640, N2384, N5148);
nand NAND2_290 (N704, N2831, N5382);
nand NAND2_291 (N1024, N3278, N2350);
nand NAND2_292 (N1216, N3427, N2585);
nand NAND2_293 (N1408, N1500, N3760);
nand NAND2_294 (N1472, N1650, N4465);
nand NAND2_295 (N650, N2400, N5170);
nand NAND2_296 (N715, N2850, N5405);
nand NAND2_297 (N1040, N3300, N2360);
nand NAND2_298 (N1235, N3450, N2596);
nand NAND2_299 (N1430, N1510, N3776);
nand NAND2_300 (N1495, N1661, N4484);
nand NAND2_301 (N660, N2416, N5192);
nand NAND2_302 (N726, N2869, N5428);
nand NAND2_303 (N1056, N3322, N2370);
nand NAND2_304 (N1254, N3473, N2607);
nand NAND2_305 (N1452, N1520, N3792);
nand NAND2_306 (N1518, N1672, N4503);
nand NAND2_307 (N670, N2432, N5214);
nand NAND2_308 (N737, N2888, N5451);
nand NAND2_309 (N1072, N3344, N2380);
nand NAND2_310 (N1273, N3496, N2618);
nand NAND2_311 (N1474, N1530, N3808);
nand NAND2_312 (N1541, N1683, N4522);
nand NAND2_313 (N680, N2448, N5236);
nand NAND2_314 (N748, N2907, N5474);
nand NAND2_315 (N1088, N3366, N2390);
nand NAND2_316 (N1292, N3519, N2629);
nand NAND2_317 (N1496, N1540, N3824);
nand NAND2_318 (N1564, N1694, N4541);
nand NAND2_319 (N690, N2464, N5258);
nand NAND2_320 (N759, N2926, N5497);
nand NAND2_321 (N1104, N3388, N2400);
nand NAND2_322 (N1311, N3542, N2640);
nand NAND2_323 (N1518, N1550, N3840);
nand NAND2_324 (N1587, N1705, N4560);
nand NAND2_325 (N700, N2480, N5280);
nand NAND2_326 (N770, N2945, N5520);
nand NAND2_327 (N1120, N3410, N2410);
nand NAND2_328 (N1330, N3565, N2651);
nand NAND2_329 (N1540, N1560, N3856);
nand NAND2_330 (N1610, N1716, N4579);
nand NAND2_331 (N710, N2496, N5302);
nand NAND2_332 (N781, N2964, N5543);
nand NAND2_333 (N1136, N3432, N2420);
nand NAND2_334 (N1349, N3588, N2662);
nand NAND2_335 (N1562, N1570, N3872);
nand NAND2_336 (N1633, N1727, N4598);
nand NAND2_337 (N720, N2512, N5324);
nand NAND2_338 (N792, N2983, N5566);
nand NAND2_339 (N1152, N3454, N2430);
nand NAND2_340 (N1368, N3611, N2673);
nand NAND2_341 (N1584, N1580, N3888);
nand NAND2_342 (N1656, N1738, N4617);
nand NAND2_343 (N730, N2528, N5346);
nand NAND2_344 (N803, N3002, N5589);
nand NAND2_345 (N1168, N3476, N2440);
nand NAND2_346 (N1387, N3634, N2684);
nand NAND2_347 (N1606, N1590, N3904);
nand NAND2_348 (N1679, N1749, N4636);
nand NAND2_349 (N740, N2544, N5368);
nand NAND2_350 (N814, N3021, N5612);
nand NAND2_351 (N1184, N3498, N2450);
nand NAND2_352 (N1406, N3657, N2695);
nand NAND2_353 (N1628, N1600, N3920);
nand NAND2_354 (N1702, N1760, N4655);
nand NAND2_355 (N750, N2560, N5390);
nand NAND2_356 (N825, N3040, N5635);
nand NAND2_357 (N1200, N3520, N2460);
nand NAND2_358 (N1425, N3680, N2706);
nand NAND2_359 (N1650, N1610, N3936);
nand NAND2_360 (N1725, N1771, N4674);
nand NAND2_361 (N760, N2576, N5412);
nand NAND2_362 (N836, N3059, N5658);
nand NAND2_363 (N1216, N3542, N2470);
nand NAND2_364 (N1444, N3703, N2717);
nand NAND2_365 (N1672, N1620, N3952);
nand NAND2_366 (N1748, N1782, N4693);
nand NAND2_367 (N770, N2592, N5434);
nand NAND2_368 (N847, N3078, N5681);
nand NAND2_369 (N1232, N3564, N2480);
nand NAND2_370 (N1463, N3726, N2728);
nand NAND2_371 (N1694, N1630, N3968);
nand NAND2_372 (N1771, N1793, N4712);
nand NAND2_373 (N780, N2608, N5456);
nand NAND2_374 (N858, N3097, N5704);
nand NAND2_375 (N1248, N3586, N2490);
nand NAND2_376 (N1482, N3749, N2739);
nand NAND2_377 (N1716, N1640, N3984);
nand NAND2_378 (N1794, N1804, N4731);
nand NAND2_379 (N790, N2624, N5478);
nand NAND2_380 (N869, N3116, N5727);
nand NAND2_381 (N1264, N3608, N2500);
nand NAND2_382 (N1501, N3772, N2750);
nand NAND2_383 (N1738, N1650, N4000);
nand NAND2_384 (N1817, N1815, N4750);
nand NAND2_385 (N800, N2640, N5500);
nand NAND2_386 (N880, N3135, N5750);
nand NAND2_387 (N1280, N3630, N2510);
nand NAND2_388 (N1520, N3795, N2761);
nand NAND2_389 (N1760, N1660, N4016);
nand NAND2_390 (N1840, N1826, N4769);
nand NAND2_391 (N810, N2656, N5522);
nand NAND2_392 (N891, N3154, N5773);
nand NAND2_393 (N1296, N3652, N2520);
nand NAND2_394 (N1539, N3818, N2772);
nand NAND2_395 (N1782, N1670, N4032);
nand NAND2_396 (N1863, N1837, N4788);
nand NAND2_397 (N820, N2672, N5544);
nand NAND2_398 (N902, N3173, N5796);
nand NAND2_399 (N1312, N3674, N2530);
nand NAND2_400 (N1558, N3841, N2783);
nand NAND2_401 (N1804, N1680, N4048);
nand NAND2_402 (N1886, N1848, N4807);
nand NAND2_403 (N830, N2688, N5566);
nand NAND2_404 (N913, N3192, N5819);
nand NAND2_405 (N1328, N3696, N2540);
nand NAND2_406 (N1577, N3864, N2794);
nand NAND2_407 (N1826, N1690, N4064);
nand NAND2_408 (N1909, N1859, N4826);
nand NAND2_409 (N840, N2704, N5588);
nand NAND2_410 (N924, N3211, N5842);
nand NAND2_411 (N1344, N3718, N2550);
nand NAND2_412 (N1596, N3887, N2805);
nand NAND2_413 (N1848, N1700, N4080);
nand NAND2_414 (N1932, N1870, N4845);
nand NAND2_415 (N850, N2720, N5610);
nand NAND2_416 (N935, N3230, N5865);
nand NAND2_417 (N1360, N3740, N2560);
nand NAND2_418 (N1615, N3910, N2816);
nand NAND2_419 (N1870, N1710, N4096);
nand NAND2_420 (N1955, N1881, N4864);
nand NAND2_421 (N860, N2736, N5632);
nand NAND2_422 (N946, N3249, N5888);
nand NAND2_423 (N1376, N3762, N2570);
nand NAND2_424 (N1634, N3933, N2827);
nand NAND2_425 (N1892, N1720, N4112);
nand NAND2_426 (N1978, N1892, N4883);
nand NAND2_427 (N870, N2752, N5654);
nand NAND2_428 (N957, N3268, N5911);
nand NAND2_429 (N1392, N3784, N2580);
nand NAND2_430 (N1653, N3956, N2838);
nand NAND2_431 (N1914, N1730, N4128);
nand NAND2_432 (N2001, N1903, N4902);
nand NAND2_433 (N880, N2768, N5676);
nand NAND2_434 (N968, N3287, N5934);
nand NAND2_435 (N1408, N3806, N2590);
nand NAND2_436 (N1672, N3979, N2849);
nand NAND2_437 (N1936, N1740, N4144);
nand NAND2_438 (N2024, N1914, N4921);
nand NAND2_439 (N890, N2784, N5698);
nand NAND2_440 (N979, N3306, N5957);
nand NAND2_441 (N1424, N3828, N2600);
nand NAND2_442 (N1691, N4002, N2860);
nand NAND2_443 (N1958, N1750, N4160);
nand NAND2_444 (N2047, N1925, N4940);
nand NAND2_445 (N900, N2800, N5720);
nand NAND2_446 (N990, N3325, N5980);
nand NAND2_447 (N1440, N3850, N2610);
nand NAND2_448 (N1710, N4025, N2871);
nand NAND2_449 (N1980, N1760, N4176);
nand NAND2_450 (N2070, N1936, N4959);
nand NAND2_451 (N910, N2816, N5742);
nand NAND2_452 (N1001, N3344, N6003);
nand NAND2_453 (N1456, N3872, N2620);
nand NAND2_454 (N1729, N4048, N2882);
nand NAND2_455 (N2002, N1770, N4192);
nand NAND2_456 (N2093, N1947, N4978);
nand NAND2_457 (N920, N2832, N5764);
nand NAND2_458 (N1012, N3363, N6026);
nand NAND2_459 (N1472, N3894, N2630);
nand NAND2_460 (N1748, N4071, N2893);
nand NAND2_461 (N2024, N1780, N4208);
nand NAND2_462 (N2116, N1958, N4997);
nand NAND2_463 (N930, N2848, N5786);
nand NAND2_464 (N1023, N3382, N6049);
nand NAND2_465 (N1488, N3916, N2640);
nand NAND2_466 (N1767, N4094, N2904);
nand NAND2_467 (N2046, N1790, N4224);
nand NAND2_468 (N2139, N1969, N5016);
nand NAND2_469 (N940, N2864, N5808);
nand NAND2_470 (N1034, N3401, N6072);
nand NAND2_471 (N1504, N3938, N2650);
nand NAND2_472 (N1786, N4117, N2915);
nand NAND2_473 (N2068, N1800, N4240);
nand NAND2_474 (N2162, N1980, N5035);
nand NAND2_475 (N950, N2880, N5830);
nand NAND2_476 (N1045, N3420, N6095);
nand NAND2_477 (N1520, N3960, N1800);
nand NAND2_478 (N1805, N4140, N2880);
nand NAND2_479 (N2090, N1810, N181);
nand NAND2_480 (N2185, N1991, N543);
nand NAND2_481 (N960, N2896, N362);
nand NAND2_482 (N1056, N3439, N1991);
nand NAND2_483 (N1536, N3982, N1810);
nand NAND2_484 (N1824, N4163, N2896);
nand NAND2_485 (N2112, N1820, N182);
nand NAND2_486 (N2208, N2002, N546);
nand NAND2_487 (N970, N2912, N364);
nand NAND2_488 (N1067, N3458, N2002);
nand NAND2_489 (N1552, N4004, N1820);
nand NAND2_490 (N1843, N4186, N2912);
nand NAND2_491 (N2134, N1830, N183);
nand NAND2_492 (N2231, N2013, N549);
nand NAND2_493 (N980, N2928, N366);
nand NAND2_494 (N1078, N3477, N2013);
nand NAND2_495 (N1568, N4026, N1830);
nand NAND2_496 (N1862, N4209, N2928);
nand NAND2_497 (N2156, N1840, N184);
nand NAND2_498 (N2254, N2024, N552);
nand NAND2_499 (N990, N2944, N368);
nand NAND2_500 (N1089, N3496, N2024);
nand NAND2_501 (N1584, N4048, N1840);
nand NAND2_502 (N1881, N4232, N2944);
nand NAND2_503 (N2178, N1850, N185);
nand NAND2_504 (N2277, N2035, N555);
nand NAND2_505 (N1000, N2960, N370);
nand NAND2_506 (N1100, N3515, N2035);
nand NAND2_507 (N1600, N4070, N1850);
nand NAND2_508 (N1900, N4255, N2960);
nand NAND2_509 (N2200, N1860, N186);
nand NAND2_510 (N2300, N2046, N558);
nand NAND2_511 (N1010, N2976, N372);
nand NAND2_512 (N1111, N3534, N2046);
nand NAND2_513 (N1616, N4092, N1860);
nand NAND2_514 (N1919, N4278, N2976);
nand NAND2_515 (N2222, N1870, N187);
nand NAND2_516 (N2323, N2057, N561);
nand NAND2_517 (N1020, N2992, N374);
nand NAND2_518 (N1122, N3553, N2057);
nand NAND2_519 (N1632, N4114, N1870);
nand NAND2_520 (N1938, N4301, N2992);
nand NAND2_521 (N2244, N1880, N188);
nand NAND2_522 (N2346, N2068, N564);
nand NAND2_523 (N1030, N3008, N376);
nand NAND2_524 (N1133, N3572, N2068);
nand NAND2_525 (N1648, N4136, N1880);
nand NAND2_526 (N1957, N4324, N3008);
nand NAND2_527 (N2266, N1890, N189);
nand NAND2_528 (N2369, N2079, N567);
nand NAND2_529 (N1040, N3024, N378);
nand NAND2_530 (N1144, N3591, N2079);
nand NAND2_531 (N1664, N4158, N1890);
nand NAND2_532 (N1976, N4347, N3024);
nand NAND2_533 (N2288, N1900, N190);
nand NAND2_534 (N2392, N2090, N570);
nand NAND2_535 (N1050, N3040, N380);
nand NAND2_536 (N1155, N3610, N2090);
nand NAND2_537 (N1680, N4180, N1900);
nand NAND2_538 (N1995, N4370, N3040);
nand NAND2_539 (N2310, N1910, N191);
nand NAND2_540 (N2415, N2101, N573);
nand NAND2_541 (N1060, N3056, N382);
nand NAND2_542 (N1166, N3629, N2101);
nand NAND2_543 (N1696, N4202, N1910);
nand NAND2_544 (N2014, N4393, N3056);
nand NAND2_545 (N2332, N1920, N192);
nand NAND2_546 (N2438, N2112, N576);
nand NAND2_547 (N1070, N3072, N384);
nand NAND2_548 (N1177, N3648, N2112);
nand NAND2_549 (N1712, N4224, N1920);
nand NAND2_550 (N2033, N4416, N3072);
nand NAND2_551 (N2354, N1930, N193);
nand NAND2_552 (N2461, N2123, N579);
nand NAND2_553 (N1080, N3088, N386);
nand NAND2_554 (N1188, N3667, N2123);
nand NAND2_555 (N1728, N4246, N1930);
nand NAND2_556 (N2052, N4439, N3088);
nand NAND2_557 (N2376, N1940, N194);
nand NAND2_558 (N2484, N2134, N582);
nand NAND2_559 (N1090, N3104, N388);
nand NAND2_560 (N1199, N3686, N2134);
nand NAND2_561 (N1744, N4268, N1940);
nand NAND2_562 (N2071, N4462, N3104);
nand NAND2_563 (N2398, N1950, N195);
nand NAND2_564 (N2507, N2145, N585);
nand NAND2_565 (N1100, N3120, N390);
nand NAND2_566 (N1210, N3705, N2145);
nand NAND2_567 (N1760, N4290, N1950);
nand NAND2_568 (N2090, N4485, N3120);
nand NAND2_569 (N2420, N1960, N196);
nand NAND2_570 (N2530, N2156, N588);
nand NAND2_571 (N1110, N3136, N392);
nand NAND2_572 (N1221, N3724, N2156);
nand NAND2_573 (N1776, N4312, N1960);
nand NAND2_574 (N2109, N4508, N3136);
nand NAND2_575 (N2442, N1970, N197);
nand NAND2_576 (N2553, N2167, N591);
nand NAND2_577 (N1120, N3152, N394);
nand NAND2_578 (N1232, N3743, N2167);
nand NAND2_579 (N1792, N4334, N1970);
nand NAND2_580 (N2128, N4531, N3152);
nand NAND2_581 (N2464, N1980, N198);
nand NAND2_582 (N2576, N2178, N594);
nand NAND2_583 (N1130, N3168, N396);
nand NAND2_584 (N1243, N3762, N2178);
nand NAND2_585 (N1808, N4356, N1980);
nand NAND2_586 (N2147, N4554, N3168);
nand NAND2_587 (N2486, N1990, N199);
nand NAND2_588 (N2599, N2189, N597);
nand NAND2_589 (N1140, N3184, N398);
nand NAND2_590 (N1254, N3781, N2189);
nand NAND2_591 (N1824, N4378, N1990);
nand NAND2_592 (N2166, N4577, N3184);
nand NAND2_593 (N2508, N2000, N200);
nand NAND2_594 (N2622, N2200, N600);
nand NAND2_595 (N1150, N3200, N400);
nand NAND2_596 (N1265, N3800, N2200);
nand NAND2_597 (N1840, N4400, N2000);
nand NAND2_598 (N2185, N4600, N3200);
nand NAND2_599 (N2530, N2010, N201);
nand NAND2_600 (N2645, N2211, N603);
nand NAND2_601 (N1160, N3216, N402);
nand NAND2_602 (N1276, N3819, N2211);
nand NAND2_603 (N1856, N4422, N2010);
nand NAND2_604 (N2204, N4623, N3216);
nand NAND2_605 (N2552, N2020, N202);
nand NAND2_606 (N2668, N2222, N606);
nand NAND2_607 (N1170, N3232, N404);
nand NAND2_608 (N1287, N3838, N2222);
nand NAND2_609 (N1872, N4444, N2020);
nand NAND2_610 (N2223, N4646, N3232);
nand NAND2_611 (N2574, N2030, N203);
nand NAND2_612 (N2691, N2233, N609);
nand NAND2_613 (N1180, N3248, N406);
nand NAND2_614 (N1298, N3857, N2233);
nand NAND2_615 (N1888, N4466, N2030);
nand NAND2_616 (N2242, N4669, N3248);
nand NAND2_617 (N2596, N2040, N204);
nand NAND2_618 (N2714, N2244, N612);
nand NAND2_619 (N1190, N3264, N408);
nand NAND2_620 (N1309, N3876, N2244);
nand NAND2_621 (N1904, N4488, N2040);
nand NAND2_622 (N2261, N4692, N3264);
nand NAND2_623 (N2618, N2050, N205);
nand NAND2_624 (N2737, N2255, N615);
nand NAND2_625 (N1200, N3280, N410);
nand NAND2_626 (N1320, N3895, N2255);
nand NAND2_627 (N1920, N4510, N2050);
nand NAND2_628 (N2280, N4715, N3280);
nand NAND2_629 (N2640, N2060, N206);
nand NAND2_630 (N2760, N2266, N618);
nand NAND2_631 (N1210, N3296, N412);
nand NAND2_632 (N1331, N3914, N2266);
nand NAND2_633 (N1936, N4532, N2060);
nand NAND2_634 (N2299, N4738, N3296);
nand NAND2_635 (N2662, N2070, N207);
nand NAND2_636 (N2783, N2277, N621);
nand NAND2_637 (N1220, N3312, N414);
nand NAND2_638 (N1342, N3933, N2277);
nand NAND2_639 (N1952, N4554, N2070);
nand NAND2_640 (N2318, N4761, N3312);
nand NAND2_641 (N2684, N2080, N208);
nand NAND2_642 (N2806, N2288, N624);
nand NAND2_643 (N1230, N3328, N416);
nand NAND2_644 (N1353, N3952, N2288);
nand NAND2_645 (N1968, N4576, N2080);
nand NAND2_646 (N2337, N4784, N3328);
nand NAND2_647 (N2706, N2090, N209);
nand NAND2_648 (N2829, N2299, N627);
nand NAND2_649 (N1240, N3344, N418);
nand NAND2_650 (N1364, N3971, N2299);
nand NAND2_651 (N1984, N4598, N2090);
nand NAND2_652 (N2356, N4807, N3344);
nand NAND2_653 (N2728, N2100, N210);
nand NAND2_654 (N2852, N2310, N630);
nand NAND2_655 (N1250, N3360, N420);
nand NAND2_656 (N1375, N3990, N2310);
nand NAND2_657 (N2000, N4620, N2100);
nand NAND2_658 (N2375, N4830, N3360);
nand NAND2_659 (N2750, N2110, N211);
nand NAND2_660 (N2875, N2321, N633);
nand NAND2_661 (N1260, N3376, N422);
nand NAND2_662 (N1386, N4009, N2321);
nand NAND2_663 (N2016, N4642, N2110);
nand NAND2_664 (N2394, N4853, N3376);
nand NAND2_665 (N2772, N2120, N212);
nand NAND2_666 (N2898, N2332, N636);
nand NAND2_667 (N1270, N3392, N424);
nand NAND2_668 (N1397, N4028, N2332);
nand NAND2_669 (N2032, N4664, N2120);
nand NAND2_670 (N2413, N4876, N3392);
nand NAND2_671 (N2794, N2130, N213);
nand NAND2_672 (N2921, N2343, N639);
nand NAND2_673 (N1280, N3408, N426);
nand NAND2_674 (N1408, N4047, N2343);
nand NAND2_675 (N2048, N4686, N2130);
nand NAND2_676 (N2432, N4899, N3408);
nand NAND2_677 (N2816, N2140, N214);
nand NAND2_678 (N2944, N2354, N642);
nand NAND2_679 (N1290, N3424, N428);
nand NAND2_680 (N1419, N4066, N2354);
nand NAND2_681 (N2064, N4708, N2140);
nand NAND2_682 (N2451, N4922, N3424);
nand NAND2_683 (N2838, N2150, N215);
nand NAND2_684 (N2967, N2365, N645);
nand NAND2_685 (N1300, N3440, N430);
nand NAND2_686 (N1430, N4085, N2365);
nand NAND2_687 (N2080, N4730, N2150);
nand NAND2_688 (N2470, N4945, N3440);
nand NAND2_689 (N2860, N2160, N216);
nand NAND2_690 (N2990, N2376, N648);
nand NAND2_691 (N1310, N3456, N432);
nand NAND2_692 (N1441, N4104, N2376);
nand NAND2_693 (N2096, N4752, N2160);
nand NAND2_694 (N2489, N4968, N3456);
nand NAND2_695 (N2882, N2170, N217);
nand NAND2_696 (N3013, N2387, N651);
nand NAND2_697 (N1320, N3472, N434);
nand NAND2_698 (N1452, N4123, N2387);
nand NAND2_699 (N2112, N4774, N2170);
nand NAND2_700 (N2508, N4991, N3472);
nand NAND2_701 (N2904, N2180, N218);
nand NAND2_702 (N3036, N2398, N654);
nand NAND2_703 (N1330, N3488, N436);
nand NAND2_704 (N1463, N4142, N2398);
nand NAND2_705 (N2128, N4796, N2180);
nand NAND2_706 (N2527, N5014, N3488);
nand NAND2_707 (N2926, N2190, N219);
nand NAND2_708 (N3059, N2409, N657);
nand NAND2_709 (N1340, N3504, N438);
nand NAND2_710 (N1474, N4161, N2409);
nand NAND2_711 (N2144, N4818, N2190);
nand NAND2_712 (N2546, N5037, N3504);
nand NAND2_713 (N2948, N2200, N220);
nand NAND2_714 (N3082, N2420, N660);
nand NAND2_715 (N1350, N3520, N440);
nand NAND2_716 (N1485, N4180, N2420);
nand NAND2_717 (N2160, N4840, N2200);
nand NAND2_718 (N2565, N5060, N3520);
nand NAND2_719 (N2970, N2210, N221);
nand NAND2_720 (N3105, N2431, N663);
nand NAND2_721 (N1360, N3536, N442);
nand NAND2_722 (N1496, N4199, N2431);
nand NAND2_723 (N2176, N4862, N2210);
nand NAND2_724 (N2584, N5083, N3536);
nand NAND2_725 (N2992, N2220, N222);
nand NAND2_726 (N3128, N2442, N666);
nand NAND2_727 (N1370, N3552, N444);
nand NAND2_728 (N1507, N4218, N2442);
nand NAND2_729 (N2192, N4884, N2220);
nand NAND2_730 (N2603, N5106, N3552);
nand NAND2_731 (N3014, N2230, N223);
nand NAND2_732 (N3151, N2453, N669);
nand NAND2_733 (N1380, N3568, N446);
nand NAND2_734 (N1518, N4237, N2453);
nand NAND2_735 (N2208, N4906, N2230);
nand NAND2_736 (N2622, N5129, N3568);
nand NAND2_737 (N3036, N2240, N224);
nand NAND2_738 (N3174, N2464, N672);
nand NAND2_739 (N1390, N3584, N448);
nand NAND2_740 (N1529, N4256, N2464);
nand NAND2_741 (N2224, N4928, N2240);
nand NAND2_742 (N2641, N5152, N3584);
nand NAND2_743 (N3058, N2250, N225);
nand NAND2_744 (N3197, N2475, N675);
nand NAND2_745 (N1400, N3600, N450);
nand NAND2_746 (N1540, N4275, N2475);
nand NAND2_747 (N2240, N4950, N2250);
nand NAND2_748 (N2660, N5175, N3600);
nand NAND2_749 (N3080, N2260, N226);
nand NAND2_750 (N3220, N2486, N678);
nand NAND2_751 (N1410, N3616, N452);
nand NAND2_752 (N1551, N4294, N2486);
nand NAND2_753 (N2256, N4972, N2260);
nand NAND2_754 (N2679, N5198, N3616);
nand NAND2_755 (N3102, N2270, N227);
nand NAND2_756 (N3243, N2497, N681);
nand NAND2_757 (N1420, N3632, N454);
nand NAND2_758 (N1562, N4313, N2497);
nand NAND2_759 (N2272, N4994, N2270);
nand NAND2_760 (N2698, N5221, N3632);
nand NAND2_761 (N3124, N2280, N228);
nand NAND2_762 (N3266, N2508, N684);
nand NAND2_763 (N1430, N3648, N456);
nand NAND2_764 (N1573, N4332, N2508);
nand NAND2_765 (N2288, N5016, N2280);
nand NAND2_766 (N2717, N5244, N3648);
nand NAND2_767 (N3146, N2290, N229);
nand NAND2_768 (N3289, N2519, N687);
nand NAND2_769 (N1440, N3664, N458);
nand NAND2_770 (N1584, N4351, N2519);
nand NAND2_771 (N2304, N5038, N2290);
nand NAND2_772 (N2736, N5267, N3664);
nand NAND2_773 (N3168, N2300, N230);
nand NAND2_774 (N3312, N2530, N690);
nand NAND2_775 (N1450, N3680, N460);
nand NAND2_776 (N1595, N4370, N2530);
nand NAND2_777 (N2320, N5060, N2300);
nand NAND2_778 (N2755, N5290, N3680);
nand NAND2_779 (N3190, N2310, N231);
nand NAND2_780 (N3335, N2541, N693);
nand NAND2_781 (N1460, N3696, N462);
nand NAND2_782 (N1606, N4389, N2541);
nand NAND2_783 (N2336, N5082, N2310);
nand NAND2_784 (N2774, N5313, N3696);
nand NAND2_785 (N3212, N2320, N232);
nand NAND2_786 (N3358, N2552, N696);
nand NAND2_787 (N1470, N3712, N464);
nand NAND2_788 (N1617, N4408, N2552);
nand NAND2_789 (N2352, N5104, N2320);
nand NAND2_790 (N2793, N5336, N3712);
nand NAND2_791 (N3234, N2330, N233);
nand NAND2_792 (N3381, N2563, N699);
nand NAND2_793 (N1480, N3728, N466);
nand NAND2_794 (N1628, N4427, N2563);
nand NAND2_795 (N2368, N5126, N2330);
nand NAND2_796 (N2812, N5359, N3728);
nand NAND2_797 (N3256, N2340, N234);
nand NAND2_798 (N3404, N2574, N702);
nand NAND2_799 (N1490, N3744, N468);
nand NAND2_800 (N1639, N4446, N2574);
nand NAND2_801 (N2384, N5148, N2340);
nand NAND2_802 (N2831, N5382, N3744);
nand NAND2_803 (N3278, N2350, N235);
nand NAND2_804 (N3427, N2585, N705);
nand NAND2_805 (N1500, N3760, N470);
nand NAND2_806 (N1650, N4465, N2585);
nand NAND2_807 (N2400, N5170, N2350);
nand NAND2_808 (N2850, N5405, N3760);
nand NAND2_809 (N3300, N2360, N236);
nand NAND2_810 (N3450, N2596, N708);
nand NAND2_811 (N1510, N3776, N472);
nand NAND2_812 (N1661, N4484, N2596);
nand NAND2_813 (N2416, N5192, N2360);
nand NAND2_814 (N2869, N5428, N3776);
nand NAND2_815 (N3322, N2370, N237);
nand NAND2_816 (N3473, N2607, N711);
nand NAND2_817 (N1520, N3792, N474);
nand NAND2_818 (N1672, N4503, N2607);
nand NAND2_819 (N2432, N5214, N2370);
nand NAND2_820 (N2888, N5451, N3792);
nand NAND2_821 (N3344, N2380, N238);
nand NAND2_822 (N3496, N2618, N714);
nand NAND2_823 (N1530, N3808, N476);
nand NAND2_824 (N1683, N4522, N2618);
nand NAND2_825 (N2448, N5236, N2380);
nand NAND2_826 (N2907, N5474, N3808);
nand NAND2_827 (N3366, N2390, N239);
nand NAND2_828 (N3519, N2629, N717);
nand NAND2_829 (N1540, N3824, N478);
nand NAND2_830 (N1694, N4541, N2629);
nand NAND2_831 (N2464, N5258, N2390);
nand NAND2_832 (N2926, N5497, N3824);
nand NAND2_833 (N3388, N2400, N240);
nand NAND2_834 (N3542, N2640, N720);
nand NAND2_835 (N1550, N3840, N480);
nand NAND2_836 (N1705, N4560, N2640);
nand NAND2_837 (N2480, N5280, N2400);
nand NAND2_838 (N2945, N5520, N3840);
nand NAND2_839 (N3410, N2410, N241);
nand NAND2_840 (N3565, N2651, N723);
nand NAND2_841 (N1560, N3856, N482);
nand NAND2_842 (N1716, N4579, N2651);
nand NAND2_843 (N2496, N5302, N2410);
nand NAND2_844 (N2964, N5543, N3856);
nand NAND2_845 (N3432, N2420, N242);
nand NAND2_846 (N3588, N2662, N726);
nand NAND2_847 (N1570, N3872, N484);
nand NAND2_848 (N1727, N4598, N2662);
nand NAND2_849 (N2512, N5324, N2420);
nand NAND2_850 (N2983, N5566, N3872);
nand NAND2_851 (N3454, N2430, N243);
nand NAND2_852 (N3611, N2673, N729);
nand NAND2_853 (N1580, N3888, N486);
nand NAND2_854 (N1738, N4617, N2673);
nand NAND2_855 (N2528, N5346, N2430);
nand NAND2_856 (N3002, N5589, N3888);
nand NAND2_857 (N3476, N2440, N244);
nand NAND2_858 (N3634, N2684, N732);
nand NAND2_859 (N1590, N3904, N488);
nand NAND2_860 (N1749, N4636, N2684);
nand NAND2_861 (N2544, N5368, N2440);
nand NAND2_862 (N3021, N5612, N3904);
nand NAND2_863 (N3498, N2450, N245);
nand NAND2_864 (N3657, N2695, N735);
nand NAND2_865 (N1600, N3920, N490);
nand NAND2_866 (N1760, N4655, N2695);
nand NAND2_867 (N2560, N5390, N2450);
nand NAND2_868 (N3040, N5635, N3920);
nand NAND2_869 (N3520, N2460, N246);
nand NAND2_870 (N3680, N2706, N738);
nand NAND2_871 (N1610, N3936, N492);
nand NAND2_872 (N1771, N4674, N2706);
nand NAND2_873 (N2576, N5412, N2460);
nand NAND2_874 (N3059, N5658, N3936);
nand NAND2_875 (N3542, N2470, N247);
nand NAND2_876 (N3703, N2717, N741);
nand NAND2_877 (N1620, N3952, N494);
nand NAND2_878 (N1782, N4693, N2717);
nand NAND2_879 (N2592, N5434, N2470);
nand NAND2_880 (N3078, N5681, N3952);
nand NAND2_881 (N3564, N2480, N248);
nand NAND2_882 (N3726, N2728, N744);
nand NAND2_883 (N1630, N3968, N496);
nand NAND2_884 (N1793, N4712, N2728);
nand NAND2_885 (N2608, N5456, N2480);
nand NAND2_886 (N3097, N5704, N3968);
nand NAND2_887 (N3586, N2490, N249);
nand NAND2_888 (N3749, N2739, N747);
nand NAND2_889 (N1640, N3984, N498);
nand NAND2_890 (N1804, N4731, N2739);
nand NAND2_891 (N2624, N5478, N2490);
nand NAND2_892 (N3116, N5727, N3984);
nand NAND2_893 (N3608, N2500, N250);
nand NAND2_894 (N3772, N2750, N750);
nand NAND2_895 (N1650, N4000, N500);
nand NAND2_896 (N1815, N4750, N2750);
nand NAND2_897 (N2640, N5500, N2500);
nand NAND2_898 (N3135, N5750, N4000);
nand NAND2_899 (N3630, N2510, N251);
nand NAND2_900 (N3795, N2761, N753);
nand NAND2_901 (N1660, N4016, N502);
nand NAND2_902 (N1826, N4769, N2761);
nand NAND2_903 (N2656, N5522, N2510);
nand NAND2_904 (N3154, N5773, N4016);
nand NAND2_905 (N3652, N2520, N252);
nand NAND2_906 (N3818, N2772, N756);
nand NAND2_907 (N1670, N4032, N504);
nand NAND2_908 (N1837, N4788, N2772);
nand NAND2_909 (N2672, N5544, N2520);
nand NAND2_910 (N3173, N5796, N4032);
nand NAND2_911 (N3674, N2530, N253);
nand NAND2_912 (N3841, N2783, N759);
nand NAND2_913 (N1680, N4048, N506);
nand NAND2_914 (N1848, N4807, N2783);
nand NAND2_915 (N2688, N5566, N2530);
nand NAND2_916 (N3192, N5819, N4048);
nand NAND2_917 (N3696, N2540, N254);
nand NAND2_918 (N3864, N2794, N762);
nand NAND2_919 (N1690, N4064, N508);
nand NAND2_920 (N1859, N4826, N2794);
nand NAND2_921 (N2704, N5588, N2540);
nand NAND2_922 (N3211, N5842, N4064);
nand NAND2_923 (N3718, N2550, N255);
nand NAND2_924 (N3887, N2805, N765);
nand NAND2_925 (N1700, N4080, N510);
nand NAND2_926 (N1870, N4845, N2805);
nand NAND2_927 (N2720, N5610, N2550);
nand NAND2_928 (N3230, N5865, N4080);
nand NAND2_929 (N3740, N2560, N256);
nand NAND2_930 (N3910, N2816, N768);
nand NAND2_931 (N1710, N4096, N512);
nand NAND2_932 (N1881, N4864, N2816);
nand NAND2_933 (N2736, N5632, N2560);
nand NAND2_934 (N3249, N5888, N4096);
nand NAND2_935 (N3762, N2570, N257);
nand NAND2_936 (N3933, N2827, N771);
nand NAND2_937 (N1720, N4112, N514);
nand NAND2_938 (N1892, N4883, N2827);
nand NAND2_939 (N2752, N5654, N2570);
nand NAND2_940 (N3268, N5911, N4112);
nand NAND2_941 (N3784, N2580, N258);
nand NAND2_942 (N3956, N2838, N774);
nand NAND2_943 (N1730, N4128, N516);
nand NAND2_944 (N1903, N4902, N2838);
nand NAND2_945 (N2768, N5676, N2580);
nand NAND2_946 (N3287, N5934, N4128);
nand NAND2_947 (N3806, N2590, N259);
nand NAND2_948 (N3979, N2849, N777);
nand NAND2_949 (N1740, N4144, N518);
nand NAND2_950 (N1914, N4921, N2849);
nand NAND2_951 (N2784, N5698, N2590);
nand NAND2_952 (N3306, N5957, N4144);
nand NAND2_953 (N3828, N2600, N260);
nand NAND2_954 (N4002, N2860, N780);
nand NAND2_955 (N1750, N4160, N520);
nand NAND2_956 (N1925, N4940, N2860);
nand NAND2_957 (N2800, N5720, N2600);
nand NAND2_958 (N3325, N5980, N4160);
nand NAND2_959 (N3850, N2610, N261);
nand NAND2_960 (N4025, N2871, N783);
nand NAND2_961 (N1760, N4176, N522);
nand NAND2_962 (N1936, N4959, N2871);
nand NAND2_963 (N2816, N5742, N2610);
nand NAND2_964 (N3344, N6003, N4176);
nand NAND2_965 (N3872, N2620, N262);
nand NAND2_966 (N4048, N2882, N786);
nand NAND2_967 (N1770, N4192, N524);
nand NAND2_968 (N1947, N4978, N2882);
nand NAND2_969 (N2832, N5764, N2620);
nand NAND2_970 (N3363, N6026, N4192);
nand NAND2_971 (N3894, N2630, N263);
nand NAND2_972 (N4071, N2893, N789);
nand NAND2_973 (N1780, N4208, N526);
nand NAND2_974 (N1958, N4997, N2893);
nand NAND2_975 (N2848, N5786, N2630);
nand NAND2_976 (N3382, N6049, N4208);
nand NAND2_977 (N3916, N2640, N264);
nand NAND2_978 (N4094, N2904, N792);
nand NAND2_979 (N1790, N4224, N528);
nand NAND2_980 (N1969, N5016, N2904);
nand NAND2_981 (N2864, N5808, N2640);
nand NAND2_982 (N3401, N6072, N4224);
nand NAND2_983 (N3938, N2650, N265);
nand NAND2_984 (N4117, N2915, N795);
nand NAND2_985 (N1800, N4240, N530);
nand NAND2_986 (N1980, N5035, N2915);
nand NAND2_987 (N2880, N5830, N2650);
nand NAND2_988 (N3420, N6095, N4240);
nand NAND2_989 (N3960, N1800, N2880);
nand NAND2_990 (N4140, N2880, N3420);
nand NAND2_991 (N1810, N181, N543);
nand NAND2_992 (N1991, N543, N1086);
nand NAND2_993 (N2896, N362, N1991);
nand NAND2_994 (N3439, N1991, N1267);
nand NAND2_995 (N3982, N1810, N2896);
nand NAND2_996 (N4163, N2896, N3439);
nand NAND2_997 (N1820, N182, N546);
nand NAND2_998 (N2002, N546, N1092);
nand NAND2_999 (N2912, N364, N2002);
nand NAND2_1000 (N3458, N2002, N1274);
nand NAND2_1001 (N4004, N1820, N2912);
nand NAND2_1002 (N4186, N2912, N3458);
nand NAND2_1003 (N1830, N183, N549);
nand NAND2_1004 (N2013, N549, N1098);
nand NAND2_1005 (N2928, N366, N2013);
nand NAND2_1006 (N3477, N2013, N1281);
nand NAND2_1007 (N4026, N1830, N2928);
nand NAND2_1008 (N4209, N2928, N3477);
nand NAND2_1009 (N1840, N184, N552);
nand NAND2_1010 (N2024, N552, N1104);
nand NAND2_1011 (N2944, N368, N2024);
nand NAND2_1012 (N3496, N2024, N1288);
nand NAND2_1013 (N4048, N1840, N2944);
nand NAND2_1014 (N4232, N2944, N3496);
nand NAND2_1015 (N1850, N185, N555);
nand NAND2_1016 (N2035, N555, N1110);
nand NAND2_1017 (N2960, N370, N2035);
nand NAND2_1018 (N3515, N2035, N1295);
nand NAND2_1019 (N4070, N1850, N2960);
nand NAND2_1020 (N4255, N2960, N3515);
nand NAND2_1021 (N1860, N186, N558);
nand NAND2_1022 (N2046, N558, N1116);
nand NAND2_1023 (N2976, N372, N2046);
nand NAND2_1024 (N3534, N2046, N1302);
nand NAND2_1025 (N4092, N1860, N2976);
nand NAND2_1026 (N4278, N2976, N3534);
nand NAND2_1027 (N1870, N187, N561);
nand NAND2_1028 (N2057, N561, N1122);
nand NAND2_1029 (N2992, N374, N2057);
nand NAND2_1030 (N3553, N2057, N1309);
nand NAND2_1031 (N4114, N1870, N2992);
nand NAND2_1032 (N4301, N2992, N3553);
nand NAND2_1033 (N1880, N188, N564);
nand NAND2_1034 (N2068, N564, N1128);
nand NAND2_1035 (N3008, N376, N2068);
nand NAND2_1036 (N3572, N2068, N1316);
nand NAND2_1037 (N4136, N1880, N3008);
nand NAND2_1038 (N4324, N3008, N3572);
nand NAND2_1039 (N1890, N189, N567);
nand NAND2_1040 (N2079, N567, N1134);
nand NAND2_1041 (N3024, N378, N2079);
nand NAND2_1042 (N3591, N2079, N1323);
nand NAND2_1043 (N4158, N1890, N3024);
nand NAND2_1044 (N4347, N3024, N3591);
nand NAND2_1045 (N1900, N190, N570);
nand NAND2_1046 (N2090, N570, N1140);
nand NAND2_1047 (N3040, N380, N2090);
nand NAND2_1048 (N3610, N2090, N1330);
nand NAND2_1049 (N4180, N1900, N3040);
nand NAND2_1050 (N4370, N3040, N3610);
nand NAND2_1051 (N1910, N191, N573);
nand NAND2_1052 (N2101, N573, N1146);
nand NAND2_1053 (N3056, N382, N2101);
nand NAND2_1054 (N3629, N2101, N1337);
nand NAND2_1055 (N4202, N1910, N3056);
nand NAND2_1056 (N4393, N3056, N3629);
nand NAND2_1057 (N1920, N192, N576);
nand NAND2_1058 (N2112, N576, N1152);
nand NAND2_1059 (N3072, N384, N2112);
nand NAND2_1060 (N3648, N2112, N1344);
nand NAND2_1061 (N4224, N1920, N3072);
nand NAND2_1062 (N4416, N3072, N3648);
nand NAND2_1063 (N1930, N193, N579);
nand NAND2_1064 (N2123, N579, N1158);
nand NAND2_1065 (N3088, N386, N2123);
nand NAND2_1066 (N3667, N2123, N1351);
nand NAND2_1067 (N4246, N1930, N3088);
nand NAND2_1068 (N4439, N3088, N3667);
nand NAND2_1069 (N1940, N194, N582);
nand NAND2_1070 (N2134, N582, N1164);
nand NAND2_1071 (N3104, N388, N2134);
nand NAND2_1072 (N3686, N2134, N1358);
nand NAND2_1073 (N4268, N1940, N3104);
nand NAND2_1074 (N4462, N3104, N3686);
nand NAND2_1075 (N1950, N195, N585);
nand NAND2_1076 (N2145, N585, N1170);
nand NAND2_1077 (N3120, N390, N2145);
nand NAND2_1078 (N3705, N2145, N1365);
nand NAND2_1079 (N4290, N1950, N3120);
nand NAND2_1080 (N4485, N3120, N3705);
nand NAND2_1081 (N1960, N196, N588);
nand NAND2_1082 (N2156, N588, N1176);
nand NAND2_1083 (N3136, N392, N2156);
nand NAND2_1084 (N3724, N2156, N1372);
nand NAND2_1085 (N4312, N1960, N3136);
nand NAND2_1086 (N4508, N3136, N3724);
nand NAND2_1087 (N1970, N197, N591);
nand NAND2_1088 (N2167, N591, N1182);
nand NAND2_1089 (N3152, N394, N2167);
nand NAND2_1090 (N3743, N2167, N1379);
nand NAND2_1091 (N4334, N1970, N3152);
nand NAND2_1092 (N4531, N3152, N3743);
nand NAND2_1093 (N1980, N198, N594);
nand NAND2_1094 (N2178, N594, N1188);
nand NAND2_1095 (N3168, N396, N2178);
nand NAND2_1096 (N3762, N2178, N1386);
nand NAND2_1097 (N4356, N1980, N3168);
nand NAND2_1098 (N4554, N3168, N3762);
nand NAND2_1099 (N1990, N199, N597);
nand NAND2_1100 (N2189, N597, N1194);
nand NAND2_1101 (N3184, N398, N2189);
nand NAND2_1102 (N3781, N2189, N1393);
nand NAND2_1103 (N4378, N1990, N3184);
nand NAND2_1104 (N4577, N3184, N3781);
nand NAND2_1105 (N2000, N200, N600);
nand NAND2_1106 (N2200, N600, N1200);
nand NAND2_1107 (N3200, N400, N2200);
nand NAND2_1108 (N3800, N2200, N1400);
nand NAND2_1109 (N4400, N2000, N3200);
nand NAND2_1110 (N4600, N3200, N3800);
nand NAND2_1111 (N2010, N201, N603);
nand NAND2_1112 (N2211, N603, N1206);
nand NAND2_1113 (N3216, N402, N2211);
nand NAND2_1114 (N3819, N2211, N1407);
nand NAND2_1115 (N4422, N2010, N3216);
nand NAND2_1116 (N4623, N3216, N3819);
nand NAND2_1117 (N2020, N202, N606);
nand NAND2_1118 (N2222, N606, N1212);
nand NAND2_1119 (N3232, N404, N2222);
nand NAND2_1120 (N3838, N2222, N1414);
nand NAND2_1121 (N4444, N2020, N3232);
nand NAND2_1122 (N4646, N3232, N3838);
nand NAND2_1123 (N2030, N203, N609);
nand NAND2_1124 (N2233, N609, N1218);
nand NAND2_1125 (N3248, N406, N2233);
nand NAND2_1126 (N3857, N2233, N1421);
nand NAND2_1127 (N4466, N2030, N3248);
nand NAND2_1128 (N4669, N3248, N3857);
nand NAND2_1129 (N2040, N204, N612);
nand NAND2_1130 (N2244, N612, N1224);
nand NAND2_1131 (N3264, N408, N2244);
nand NAND2_1132 (N3876, N2244, N1428);
nand NAND2_1133 (N4488, N2040, N3264);
nand NAND2_1134 (N4692, N3264, N3876);
nand NAND2_1135 (N2050, N205, N615);
nand NAND2_1136 (N2255, N615, N1230);
nand NAND2_1137 (N3280, N410, N2255);
nand NAND2_1138 (N3895, N2255, N1435);
nand NAND2_1139 (N4510, N2050, N3280);
nand NAND2_1140 (N4715, N3280, N3895);
nand NAND2_1141 (N2060, N206, N618);
nand NAND2_1142 (N2266, N618, N1236);
nand NAND2_1143 (N3296, N412, N2266);
nand NAND2_1144 (N3914, N2266, N1442);
nand NAND2_1145 (N4532, N2060, N3296);
nand NAND2_1146 (N4738, N3296, N3914);
nand NAND2_1147 (N2070, N207, N621);
nand NAND2_1148 (N2277, N621, N1242);
nand NAND2_1149 (N3312, N414, N2277);
nand NAND2_1150 (N3933, N2277, N1449);
nand NAND2_1151 (N4554, N2070, N3312);
nand NAND2_1152 (N4761, N3312, N3933);
nand NAND2_1153 (N2080, N208, N624);
nand NAND2_1154 (N2288, N624, N1248);
nand NAND2_1155 (N3328, N416, N2288);
nand NAND2_1156 (N3952, N2288, N1456);
nand NAND2_1157 (N4576, N2080, N3328);
nand NAND2_1158 (N4784, N3328, N3952);
nand NAND2_1159 (N2090, N209, N627);
nand NAND2_1160 (N2299, N627, N1254);
nand NAND2_1161 (N3344, N418, N2299);
nand NAND2_1162 (N3971, N2299, N1463);
nand NAND2_1163 (N4598, N2090, N3344);
nand NAND2_1164 (N4807, N3344, N3971);
nand NAND2_1165 (N2100, N210, N630);
nand NAND2_1166 (N2310, N630, N1260);
nand NAND2_1167 (N3360, N420, N2310);
nand NAND2_1168 (N3990, N2310, N1470);
nand NAND2_1169 (N4620, N2100, N3360);
nand NAND2_1170 (N4830, N3360, N3990);
nand NAND2_1171 (N2110, N211, N633);
nand NAND2_1172 (N2321, N633, N1266);
nand NAND2_1173 (N3376, N422, N2321);
nand NAND2_1174 (N4009, N2321, N1477);
nand NAND2_1175 (N4642, N2110, N3376);
nand NAND2_1176 (N4853, N3376, N4009);
nand NAND2_1177 (N2120, N212, N636);
nand NAND2_1178 (N2332, N636, N1272);
nand NAND2_1179 (N3392, N424, N2332);
nand NAND2_1180 (N4028, N2332, N1484);
nand NAND2_1181 (N4664, N2120, N3392);
nand NAND2_1182 (N4876, N3392, N4028);
nand NAND2_1183 (N2130, N213, N639);
nand NAND2_1184 (N2343, N639, N1278);
nand NAND2_1185 (N3408, N426, N2343);
nand NAND2_1186 (N4047, N2343, N1491);
nand NAND2_1187 (N4686, N2130, N3408);
nand NAND2_1188 (N4899, N3408, N4047);
nand NAND2_1189 (N2140, N214, N642);
nand NAND2_1190 (N2354, N642, N1284);
nand NAND2_1191 (N3424, N428, N2354);
nand NAND2_1192 (N4066, N2354, N1498);
nand NAND2_1193 (N4708, N2140, N3424);
nand NAND2_1194 (N4922, N3424, N4066);
nand NAND2_1195 (N2150, N215, N645);
nand NAND2_1196 (N2365, N645, N1290);
nand NAND2_1197 (N3440, N430, N2365);
nand NAND2_1198 (N4085, N2365, N1505);
nand NAND2_1199 (N4730, N2150, N3440);
nand NAND2_1200 (N4945, N3440, N4085);
nand NAND2_1201 (N2160, N216, N648);
nand NAND2_1202 (N2376, N648, N1296);
nand NAND2_1203 (N3456, N432, N2376);
nand NAND2_1204 (N4104, N2376, N1512);
nand NAND2_1205 (N4752, N2160, N3456);
nand NAND2_1206 (N4968, N3456, N4104);
nand NAND2_1207 (N2170, N217, N651);
nand NAND2_1208 (N2387, N651, N1302);
nand NAND2_1209 (N3472, N434, N2387);
nand NAND2_1210 (N4123, N2387, N1519);
nand NAND2_1211 (N4774, N2170, N3472);
nand NAND2_1212 (N4991, N3472, N4123);
nand NAND2_1213 (N2180, N218, N654);
nand NAND2_1214 (N2398, N654, N1308);
nand NAND2_1215 (N3488, N436, N2398);
nand NAND2_1216 (N4142, N2398, N1526);
nand NAND2_1217 (N4796, N2180, N3488);
nand NAND2_1218 (N5014, N3488, N4142);
nand NAND2_1219 (N2190, N219, N657);
nand NAND2_1220 (N2409, N657, N1314);
nand NAND2_1221 (N3504, N438, N2409);
nand NAND2_1222 (N4161, N2409, N1533);
nand NAND2_1223 (N4818, N2190, N3504);
nand NAND2_1224 (N5037, N3504, N4161);
nand NAND2_1225 (N2200, N220, N660);
nand NAND2_1226 (N2420, N660, N1320);
nand NAND2_1227 (N3520, N440, N2420);
nand NAND2_1228 (N4180, N2420, N1540);
nand NAND2_1229 (N4840, N2200, N3520);
nand NAND2_1230 (N5060, N3520, N4180);
nand NAND2_1231 (N2210, N221, N663);
nand NAND2_1232 (N2431, N663, N1326);
nand NAND2_1233 (N3536, N442, N2431);
nand NAND2_1234 (N4199, N2431, N1547);
nand NAND2_1235 (N4862, N2210, N3536);
nand NAND2_1236 (N5083, N3536, N4199);
nand NAND2_1237 (N2220, N222, N666);
nand NAND2_1238 (N2442, N666, N1332);
nand NAND2_1239 (N3552, N444, N2442);
nand NAND2_1240 (N4218, N2442, N1554);
nand NAND2_1241 (N4884, N2220, N3552);
nand NAND2_1242 (N5106, N3552, N4218);
nand NAND2_1243 (N2230, N223, N669);
nand NAND2_1244 (N2453, N669, N1338);
nand NAND2_1245 (N3568, N446, N2453);
nand NAND2_1246 (N4237, N2453, N1561);
nand NAND2_1247 (N4906, N2230, N3568);
nand NAND2_1248 (N5129, N3568, N4237);
nand NAND2_1249 (N2240, N224, N672);
nand NAND2_1250 (N2464, N672, N1344);
nand NAND2_1251 (N3584, N448, N2464);
nand NAND2_1252 (N4256, N2464, N1568);
nand NAND2_1253 (N4928, N2240, N3584);
nand NAND2_1254 (N5152, N3584, N4256);
nand NAND2_1255 (N2250, N225, N675);
nand NAND2_1256 (N2475, N675, N1350);
nand NAND2_1257 (N3600, N450, N2475);
nand NAND2_1258 (N4275, N2475, N1575);
nand NAND2_1259 (N4950, N2250, N3600);
nand NAND2_1260 (N5175, N3600, N4275);
nand NAND2_1261 (N2260, N226, N678);
nand NAND2_1262 (N2486, N678, N1356);
nand NAND2_1263 (N3616, N452, N2486);
nand NAND2_1264 (N4294, N2486, N1582);
nand NAND2_1265 (N4972, N2260, N3616);
nand NAND2_1266 (N5198, N3616, N4294);
nand NAND2_1267 (N2270, N227, N681);
nand NAND2_1268 (N2497, N681, N1362);
nand NAND2_1269 (N3632, N454, N2497);
nand NAND2_1270 (N4313, N2497, N1589);
nand NAND2_1271 (N4994, N2270, N3632);
nand NAND2_1272 (N5221, N3632, N4313);
nand NAND2_1273 (N2280, N228, N684);
nand NAND2_1274 (N2508, N684, N1368);
nand NAND2_1275 (N3648, N456, N2508);
nand NAND2_1276 (N4332, N2508, N1596);
nand NAND2_1277 (N5016, N2280, N3648);
nand NAND2_1278 (N5244, N3648, N4332);
nand NAND2_1279 (N2290, N229, N687);
nand NAND2_1280 (N2519, N687, N1374);
nand NAND2_1281 (N3664, N458, N2519);
nand NAND2_1282 (N4351, N2519, N1603);
nand NAND2_1283 (N5038, N2290, N3664);
nand NAND2_1284 (N5267, N3664, N4351);
nand NAND2_1285 (N2300, N230, N690);
nand NAND2_1286 (N2530, N690, N1380);
nand NAND2_1287 (N3680, N460, N2530);
nand NAND2_1288 (N4370, N2530, N1610);
nand NAND2_1289 (N5060, N2300, N3680);
nand NAND2_1290 (N5290, N3680, N4370);
nand NAND2_1291 (N2310, N231, N693);
nand NAND2_1292 (N2541, N693, N1386);
nand NAND2_1293 (N3696, N462, N2541);
nand NAND2_1294 (N4389, N2541, N1617);
nand NAND2_1295 (N5082, N2310, N3696);
nand NAND2_1296 (N5313, N3696, N4389);
nand NAND2_1297 (N2320, N232, N696);
nand NAND2_1298 (N2552, N696, N1392);
nand NAND2_1299 (N3712, N464, N2552);
nand NAND2_1300 (N4408, N2552, N1624);
nand NAND2_1301 (N5104, N2320, N3712);
nand NAND2_1302 (N5336, N3712, N4408);
nand NAND2_1303 (N2330, N233, N699);
nand NAND2_1304 (N2563, N699, N1398);
nand NAND2_1305 (N3728, N466, N2563);
nand NAND2_1306 (N4427, N2563, N1631);
nand NAND2_1307 (N5126, N2330, N3728);
nand NAND2_1308 (N5359, N3728, N4427);
nand NAND2_1309 (N2340, N234, N702);
nand NAND2_1310 (N2574, N702, N1404);
nand NAND2_1311 (N3744, N468, N2574);
nand NAND2_1312 (N4446, N2574, N1638);
nand NAND2_1313 (N5148, N2340, N3744);
nand NAND2_1314 (N5382, N3744, N4446);
nand NAND2_1315 (N2350, N235, N705);
nand NAND2_1316 (N2585, N705, N1410);
nand NAND2_1317 (N3760, N470, N2585);
nand NAND2_1318 (N4465, N2585, N1645);
nand NAND2_1319 (N5170, N2350, N3760);
nand NAND2_1320 (N5405, N3760, N4465);
nand NAND2_1321 (N2360, N236, N708);
nand NAND2_1322 (N2596, N708, N1416);
nand NAND2_1323 (N3776, N472, N2596);
nand NAND2_1324 (N4484, N2596, N1652);
nand NAND2_1325 (N5192, N2360, N3776);
nand NAND2_1326 (N5428, N3776, N4484);
nand NAND2_1327 (N2370, N237, N711);
nand NAND2_1328 (N2607, N711, N1422);
nand NAND2_1329 (N3792, N474, N2607);
nand NAND2_1330 (N4503, N2607, N1659);
nand NAND2_1331 (N5214, N2370, N3792);
nand NAND2_1332 (N5451, N3792, N4503);
nand NAND2_1333 (N2380, N238, N714);
nand NAND2_1334 (N2618, N714, N1428);
nand NAND2_1335 (N3808, N476, N2618);
nand NAND2_1336 (N4522, N2618, N1666);
nand NAND2_1337 (N5236, N2380, N3808);
nand NAND2_1338 (N5474, N3808, N4522);
nand NAND2_1339 (N2390, N239, N717);
nand NAND2_1340 (N2629, N717, N1434);
nand NAND2_1341 (N3824, N478, N2629);
nand NAND2_1342 (N4541, N2629, N1673);
nand NAND2_1343 (N5258, N2390, N3824);
nand NAND2_1344 (N5497, N3824, N4541);
nand NAND2_1345 (N2400, N240, N720);
nand NAND2_1346 (N2640, N720, N1440);
nand NAND2_1347 (N3840, N480, N2640);
nand NAND2_1348 (N4560, N2640, N1680);
nand NAND2_1349 (N5280, N2400, N3840);
nand NAND2_1350 (N5520, N3840, N4560);
nand NAND2_1351 (N2410, N241, N723);
nand NAND2_1352 (N2651, N723, N1446);
nand NAND2_1353 (N3856, N482, N2651);
nand NAND2_1354 (N4579, N2651, N1687);
nand NAND2_1355 (N5302, N2410, N3856);
nand NAND2_1356 (N5543, N3856, N4579);
nand NAND2_1357 (N2420, N242, N726);
nand NAND2_1358 (N2662, N726, N1452);
nand NAND2_1359 (N3872, N484, N2662);
nand NAND2_1360 (N4598, N2662, N1694);
nand NAND2_1361 (N5324, N2420, N3872);
nand NAND2_1362 (N5566, N3872, N4598);
nand NAND2_1363 (N2430, N243, N729);
nand NAND2_1364 (N2673, N729, N1458);
nand NAND2_1365 (N3888, N486, N2673);
nand NAND2_1366 (N4617, N2673, N1701);
nand NAND2_1367 (N5346, N2430, N3888);
nand NAND2_1368 (N5589, N3888, N4617);
nand NAND2_1369 (N2440, N244, N732);
nand NAND2_1370 (N2684, N732, N1464);
nand NAND2_1371 (N3904, N488, N2684);
nand NAND2_1372 (N4636, N2684, N1708);
nand NAND2_1373 (N5368, N2440, N3904);
nand NAND2_1374 (N5612, N3904, N4636);
nand NAND2_1375 (N2450, N245, N735);
nand NAND2_1376 (N2695, N735, N1470);
nand NAND2_1377 (N3920, N490, N2695);
nand NAND2_1378 (N4655, N2695, N1715);
nand NAND2_1379 (N5390, N2450, N3920);
nand NAND2_1380 (N5635, N3920, N4655);
nand NAND2_1381 (N2460, N246, N738);
nand NAND2_1382 (N2706, N738, N1476);
nand NAND2_1383 (N3936, N492, N2706);
nand NAND2_1384 (N4674, N2706, N1722);
nand NAND2_1385 (N5412, N2460, N3936);
nand NAND2_1386 (N5658, N3936, N4674);
nand NAND2_1387 (N2470, N247, N741);
nand NAND2_1388 (N2717, N741, N1482);
nand NAND2_1389 (N3952, N494, N2717);
nand NAND2_1390 (N4693, N2717, N1729);
nand NAND2_1391 (N5434, N2470, N3952);
nand NAND2_1392 (N5681, N3952, N4693);
nand NAND2_1393 (N2480, N248, N744);
nand NAND2_1394 (N2728, N744, N1488);
nand NAND2_1395 (N3968, N496, N2728);
nand NAND2_1396 (N4712, N2728, N1736);
nand NAND2_1397 (N5456, N2480, N3968);
nand NAND2_1398 (N5704, N3968, N4712);
nand NAND2_1399 (N2490, N249, N747);
nand NAND2_1400 (N2739, N747, N1494);
nand NAND2_1401 (N3984, N498, N2739);
nand NAND2_1402 (N4731, N2739, N1743);
nand NAND2_1403 (N5478, N2490, N3984);
nand NAND2_1404 (N5727, N3984, N4731);
nand NAND2_1405 (N2500, N250, N750);
nand NAND2_1406 (N2750, N750, N1500);
nand NAND2_1407 (N4000, N500, N2750);
nand NAND2_1408 (N4750, N2750, N1750);
nand NAND2_1409 (N5500, N2500, N4000);
nand NAND2_1410 (N5750, N4000, N4750);
nand NAND2_1411 (N2510, N251, N753);
nand NAND2_1412 (N2761, N753, N1506);
nand NAND2_1413 (N4016, N502, N2761);
nand NAND2_1414 (N4769, N2761, N1757);
nand NAND2_1415 (N5522, N2510, N4016);
nand NAND2_1416 (N5773, N4016, N4769);
nand NAND2_1417 (N2520, N252, N756);
nand NAND2_1418 (N2772, N756, N1512);
nand NAND2_1419 (N4032, N504, N2772);
nand NAND2_1420 (N4788, N2772, N1764);
nand NAND2_1421 (N5544, N2520, N4032);
nand NAND2_1422 (N5796, N4032, N4788);
nand NAND2_1423 (N2530, N253, N759);
nand NAND2_1424 (N2783, N759, N1518);
nand NAND2_1425 (N4048, N506, N2783);
nand NAND2_1426 (N4807, N2783, N1771);
nand NAND2_1427 (N5566, N2530, N4048);
nand NAND2_1428 (N5819, N4048, N4807);
nand NAND2_1429 (N2540, N254, N762);
nand NAND2_1430 (N2794, N762, N1524);
nand NAND2_1431 (N4064, N508, N2794);
nand NAND2_1432 (N4826, N2794, N1778);
nand NAND2_1433 (N5588, N2540, N4064);
nand NAND2_1434 (N5842, N4064, N4826);
nand NAND2_1435 (N2550, N255, N765);
nand NAND2_1436 (N2805, N765, N1530);
nand NAND2_1437 (N4080, N510, N2805);
nand NAND2_1438 (N4845, N2805, N1785);
nand NAND2_1439 (N5610, N2550, N4080);
nand NAND2_1440 (N5865, N4080, N4845);
nand NAND2_1441 (N2560, N256, N768);
nand NAND2_1442 (N2816, N768, N1536);
nand NAND2_1443 (N4096, N512, N2816);
nand NAND2_1444 (N4864, N2816, N1792);
nand NAND2_1445 (N5632, N2560, N4096);
nand NAND2_1446 (N5888, N4096, N4864);
nand NAND2_1447 (N2570, N257, N771);
nand NAND2_1448 (N2827, N771, N1542);
nand NAND2_1449 (N4112, N514, N2827);
nand NAND2_1450 (N4883, N2827, N1799);
nand NAND2_1451 (N5654, N2570, N4112);
nand NAND2_1452 (N5911, N4112, N4883);
nand NAND2_1453 (N2580, N258, N774);
nand NAND2_1454 (N2838, N774, N1548);
nand NAND2_1455 (N4128, N516, N2838);
nand NAND2_1456 (N4902, N2838, N1806);
nand NAND2_1457 (N5676, N2580, N4128);
nand NAND2_1458 (N5934, N4128, N4902);
nand NAND2_1459 (N2590, N259, N777);
nand NAND2_1460 (N2849, N777, N1554);
nand NAND2_1461 (N4144, N518, N2849);
nand NAND2_1462 (N4921, N2849, N1813);
nand NAND2_1463 (N5698, N2590, N4144);
nand NAND2_1464 (N5957, N4144, N4921);
nand NAND2_1465 (N2600, N260, N780);
nand NAND2_1466 (N2860, N780, N1560);
nand NAND2_1467 (N4160, N520, N2860);
nand NAND2_1468 (N4940, N2860, N1820);
nand NAND2_1469 (N5720, N2600, N4160);
nand NAND2_1470 (N5980, N4160, N4940);
nand NAND2_1471 (N2610, N261, N783);
nand NAND2_1472 (N2871, N783, N1566);
nand NAND2_1473 (N4176, N522, N2871);
nand NAND2_1474 (N4959, N2871, N1827);
nand NAND2_1475 (N5742, N2610, N4176);
nand NAND2_1476 (N6003, N4176, N4959);
nand NAND2_1477 (N2620, N262, N786);
nand NAND2_1478 (N2882, N786, N1572);
nand NAND2_1479 (N4192, N524, N2882);
nand NAND2_1480 (N4978, N2882, N1834);
nand NAND2_1481 (N5764, N2620, N4192);
nand NAND2_1482 (N6026, N4192, N4978);
nand NAND2_1483 (N2630, N263, N789);
nand NAND2_1484 (N2893, N789, N1578);
nand NAND2_1485 (N4208, N526, N2893);
nand NAND2_1486 (N4997, N2893, N1841);
nand NAND2_1487 (N5786, N2630, N4208);
nand NAND2_1488 (N6049, N4208, N4997);
nand NAND2_1489 (N2640, N264, N792);
nand NAND2_1490 (N2904, N792, N1584);
nand NAND2_1491 (N4224, N528, N2904);
nand NAND2_1492 (N5016, N2904, N1848);
nand NAND2_1493 (N5808, N2640, N4224);
nand NAND2_1494 (N6072, N4224, N5016);
nand NAND2_1495 (N2650, N265, N795);
nand NAND2_1496 (N2915, N795, N1590);
nand NAND2_1497 (N4240, N530, N2915);
nand NAND2_1498 (N5035, N2915, N1855);
nand NAND2_1499 (N5830, N2650, N4240);
nand NAND2_1500 (N6095, N4240, N5035);

endmodule
