module c34 (N1,N2,N3,N6,N7,N17,N34,N51,N102,N119,N22,N23,N374,N391);

input N1,N2,N3,N6,N7,N17,N34,N51,N102,N119;

output N22,N23,N374,N391;

wire N10,N11,N16,N19,N170,N187;

nand NAND2_1 (N10, N1, N3);
nand NAND2_2 (N11, N3, N6);
nand NAND2_3 (N16, N2, N11);
nand NAND2_4 (N19, N11, N7);
nand NAND2_5 (N22, N10, N16);
nand NAND2_6 (N23, N16, N19);
nand NAND2_7 (N170, N17, N51);
nand NAND2_8 (N187, N51, N102);
nand NAND2_9 (N272, N34, N187);
nand NAND2_10 (N323, N187, N119);
nand NAND2_11 (N374, N170, N272);
nand NAND2_12 (N391, N272, N323);

endmodule
