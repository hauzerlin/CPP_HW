module c17 (